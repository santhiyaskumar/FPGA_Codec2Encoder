/*
* Module         - ROM_cb4
* Top module     - cbselect
* Project        - CODEC2_ENCODE_2400
* Developer      - Santhiya S
* Date           - Mon Feb 04 15:19:31 2019
*
* Description    -
* Inputs         -
*static const float codes4[] = {
  950,
  1050,
  1150,
  1250,
  1350,
  1450,
  1550,
  1650,
  1750,
  1850,
  1950,
  2050,
  2150,
  2250,
  2350,
  2450
*};
*32 bits fixed point representation
   S - E  - M
   1 - 15 - 16
*/
module ROM_cb4(addr,dataout);

	parameter N = 32;
	input [3:0] addr;
	output reg [N-1:0] dataout;

	reg [N-1:0] cb4[15:0];
	
	always@(*)
	begin
		cb4[0] = 32'b00000011101101100000000000000000;
		cb4[1] = 32'b00000100000110100000000000000000;
		cb4[2] = 32'b00000100011111100000000000000000;
		cb4[3] = 32'b00000100111000100000000000000000;
		cb4[4] = 32'b00000101010001100000000000000000;
		cb4[5] = 32'b00000101101010100000000000000000;
		cb4[6] = 32'b00000110000011100000000000000000;
		cb4[7] = 32'b00000110011100100000000000000000;
		cb4[8] = 32'b00000110110101100000000000000000;
		cb4[9] = 32'b00000111001110100000000000000000;
		cb4[10] = 32'b00000111100111100000000000000000;
		cb4[11] = 32'b00001000000000100000000000000000;
		cb4[12] = 32'b00001000011001100000000000000000;
		cb4[13] = 32'b00001000110010100000000000000000;
		cb4[14] = 32'b00001001001011100000000000000000;
		cb4[15] = 32'b00001001100100100000000000000000;

		dataout = cb4[addr];
	end
endmodule
