/*
* Module         - encode_WoE
* Top module     - codec2_encode
* Project        - CODEC2_ENCODE_2400
* Developer      - Santhiya S
* Date           - Wed Feb 20 13:16:46 2019
*
* Description    -
* Inputs         -
* Simulation     - Waveform36.vwf
*32 bits fixed point representation
   S - E  - M
   1 - 15 - 16
*/


module encode_WoE (startewoe,clk,rst,model_wo,in_e,xq0,xq1,out_xq0,out_xq1,out_n1,doneewoe);
							//check_x0,check_x1,check_mult,check_logx,check_e,check_add1);


//------------------------------------------------------------------
//                 -- Input/Output Declarations --                  
//------------------------------------------------------------------

	parameter N = 32;
	parameter Q = 16;
	
	input startewoe, clk, rst;
	input [N-1:0] model_wo, in_e,xq0,xq1;
	output reg [N-1:0] out_n1,out_xq0,out_xq1;
	output reg doneewoe;
	
//	output reg [N-1:0] check_x0,check_x1,check_mult,check_logx,check_e,check_add1;

//------------------------------------------------------------------
//                  -- State & Reg Declarations  --                   
//------------------------------------------------------------------

parameter START = 5'd0,
          CHECK_E = 5'd1,
          SET_E = 5'd2,
          PRECALC1_X0 = 5'd3,
          PRECALC2_X0 = 5'd4,
          PRE_CALC3_X0 = 5'd5,
          CALC_X0 = 5'd6,
          PRECALC_X1 = 5'd7,
          CALC_X1 = 5'd8,
          SET_CW = 5'd9,
          CALC_CW = 5'd10,
          PRECALC1_ERR = 5'd11,
          PRECALC2_ERR = 5'd12,
          CALC_ERR = 5'd13,
          SET_FNW = 5'd14,
          CALC_FNW = 5'd15,
          DONE = 5'd16,
		  SET_XQ0 = 5'd17,
		  XQ0_ADD = 5'd18,
		  XQ0_MULT = 5'd19;
		  

reg [4:0]STATE, NEXT_STATE;

parameter [N-1:0] 	cb0 = 32'b00000000000000101011010111000010,
						cb1 = 32'b00000000000011000000010010110101,
						cb2 = 32'b00000000000000000000101111110111,
						cb3 = 32'b10000000000000101011110100100010,
						cb4 = 32'b00000000000000000001111011111001,
						cb5 = 32'b00000000000010000110001110010010,
						cb6 = 32'b10000000000000011001010010001101,
						cb7 = 32'b10000000000000001110010001101110,
						cb8 = 32'b00000000000000010011000101101101,
						cb9 = 32'b10000000000000011110101001100101,
						cb10 = 32'b00000000000000000010111111100101,
						cb11 = 32'b10000000000000110100011011011011,
						cb12 = 32'b00000000000000000101010100001110,
						cb13 = 32'b10000000000001111010101000011111,
						cb14 = 32'b10000000000000010111101010111100,
						cb15 = 32'b00000000000111110011111100000000,
						cb16 = 32'b00000000000000011000011100010001,
						cb17 = 32'b00000000000110111011010110100001,
						cb18 = 32'b10000000000000001000011000111101,
						cb19 = 32'b00000000000001010100000000000111,
						cb20 = 32'b00000000000000001000110110100111,
						cb21 = 32'b00000000000001110111000001010101,
						cb22 = 32'b10000000000000001101011111101100,
						cb23 = 32'b10000000000000011111001111110111,
						cb24 = 32'b00000000000000100100001110001110,
						cb25 = 32'b00000000000010001001110000111011,
						cb26 = 32'b00000000000000000010010010100101,
						cb27 = 32'b00000000000000100101110110010000,
						cb28 = 32'b00000000000000001001110111010011,
						cb29 = 32'b00000000000000010100100011000101,
						cb30 = 32'b10000000000000011011011000011001,
						cb31 = 32'b00000000000101100001100011000001,
						cb32 = 32'b00000000000000010000001000010100,
						cb33 = 32'b00000000000100010110010110000001,
						cb34 = 32'b10000000000000000001101101010001,
						cb35 = 32'b00000000000000010110101100111101,
						cb36 = 32'b10000000000000000010001011100001,
						cb37 = 32'b00000000000011100100011000001010,
						cb38 = 32'b10000000000000011011010110000110,
						cb39 = 32'b10000000000101001000100000101010,
						cb40 = 32'b00000000000000011010100001101010,
						cb41 = 32'b10000000000000110110010000011101,
						cb42 = 32'b00000000000000000010001101010111,
						cb43 = 32'b10000000000001001111010100110101,
						cb44 = 32'b00000000000000001000100101100111,
						cb45 = 32'b10000000000000011111000110011001,
						cb46 = 32'b00000000000000000011001001000001,
						cb47 = 32'b00000000001001001101101000010110,
						cb48 = 32'b00000000000000010100010111000001,
						cb49 = 32'b00000000000101101000111001110110,
						cb50 = 32'b10000000000000001010101110010011,
						cb51 = 32'b10000000000000011110011111110010,
						cb52 = 32'b00000000000000000110000111010000,
						cb53 = 32'b00000000000001100110011010110000,
						cb54 = 32'b10000000000000001100000111000100,
						cb55 = 32'b10000000000001001110011010101001,
						cb56 = 32'b00000000000000011101010001001101,
						cb57 = 32'b00000000000001001001110100100001,
						cb58 = 32'b00000000000000000101000110011100,
						cb59 = 32'b00000000000000001011110010100000,
						cb60 = 32'b00000000000000001001110011100001,
						cb61 = 32'b10000000000000100001001100110110,
						cb62 = 32'b10000000000000000110100011111111,
						cb63 = 32'b00000000000110001100100101111111,
						cb64 = 32'b00000000000000011100011010101001,
						cb65 = 32'b00000000000011010011000011011110,
						cb66 = 32'b00000000000000000001101101000000,
						cb67 = 32'b10000000000000000001101010111111,
						cb68 = 32'b00000000000000000011000100110100,
						cb69 = 32'b00000000000010100010111100001101,
						cb70 = 32'b10000000000000011101001100001101,
						cb71 = 32'b10000000000001111011011100110100,
						cb72 = 32'b00000000000000001110111001101100,
						cb73 = 32'b00000000000001000101100100101101,
						cb74 = 32'b00000000000000000100111100001110,
						cb75 = 32'b10000000000001000001011000000100,
						cb76 = 32'b00000000000000000110010110101011,
						cb77 = 32'b10000000000010111100111100010100,
						cb78 = 32'b10000000000000000000110001111000,
						cb79 = 32'b00000000001010010011101000110000,
						cb80 = 32'b00000000000000001110000010011001,
						cb81 = 32'b00000000001000111101100110101101,
						cb82 = 32'b10000000000000001100001010000001,
						cb83 = 32'b00000000000000000111101000000100,
						cb84 = 32'b00000000000000001111101010000101,
						cb85 = 32'b00000000000001111010110010110111,
						cb86 = 32'b10000000000000010011000111101111,
						cb87 = 32'b00000000000000110000100111110000,
						cb88 = 32'b00000000000000101010001111001111,
						cb89 = 32'b10000000000000110110100100111011,
						cb90 = 32'b00000000000000000011000011101101,
						cb91 = 32'b00000000000000111001101001111111,
						cb92 = 32'b00000000000000000110011100100110,
						cb93 = 32'b00000000000000010001010110010100,
						cb94 = 32'b10000000000000100010011011101010,
						cb95 = 32'b00000000000100100001101110001011,
						cb96 = 32'b00000000000000011000101111111011,
						cb97 = 32'b00000000000010000101001010011101,
						cb98 = 32'b10000000000000000010010010100001,
						cb99 = 32'b10000000000001000001001101101111,
						cb100 = 32'b10000000000000000010011001101111,
						cb101 = 32'b00000000000001011101110111100010,
						cb102 = 32'b10000000000000010110100010001111,
						cb103 = 32'b10000000000000110100000000101101,
						cb104 = 32'b00000000000000011001000011101111,
						cb105 = 32'b10000000000010100110100111000111,
						cb106 = 32'b00000000000000000010110110011100,
						cb107 = 32'b10000000000010100011101000001001,
						cb108 = 32'b00000000000000000101110010110110,
						cb109 = 32'b10000000000000000000011101001111,
						cb110 = 32'b10000000000000000001000111110011,
						cb111 = 32'b00000000000110000110010000000100,
						cb112 = 32'b00000000000000001001100001000001,
						cb113 = 32'b00000000000100010111101110011000,
						cb114 = 32'b10000000000000000100100101110111,
						cb115 = 32'b10000000000001101110011101110001,
						cb116 = 32'b00000000000000000111011011111110,
						cb117 = 32'b00000000000010100011010010011011,
						cb118 = 32'b10000000000000010000000111000000,
						cb119 = 32'b10000000000011100101101101110001,
						cb120 = 32'b00000000000000100101010001011110,
						cb121 = 32'b10000000000000111011000100001101,
						cb122 = 32'b00000000000000000101010111110011,
						cb123 = 32'b00000000000000100110100000111010,
						cb124 = 32'b00000000000000010000010100001000,
						cb125 = 32'b10000000000000110010011111011000,
						cb126 = 32'b10000000000000010100001001101011,
						cb127 = 32'b00000000000001111111110111101101,
						cb128 = 32'b00000000000000100110001000111001,
						cb129 = 32'b00000000000100111010111000111011,
						cb130 = 32'b10000000000000000001100001001110,
						cb131 = 32'b10000000000000100110100111101010,
						cb132 = 32'b00000000000000000011010110010110,
						cb133 = 32'b00000000000001101010101000101110,
						cb134 = 32'b10000000000000100011100010010101,
						cb135 = 32'b00000000000000010110000100111110,
						cb136 = 32'b00000000000000010100101011011010,
						cb137 = 32'b00000000000000100000101111011100,
						cb138 = 32'b00000000000000000011111001011110,
						cb139 = 32'b10000000000000001110010000000111,
						cb140 = 32'b00000000000000000110110111000100,
						cb141 = 32'b10000000000001110011000110010011,
						cb142 = 32'b10000000000000010001110100011110,
						cb143 = 32'b00000000001010010101011101100101,
						cb144 = 32'b00000000000000101001110000011011,
						cb145 = 32'b00000000000111110010001111110111,
						cb146 = 32'b10000000000000000111001001001011,
						cb147 = 32'b00000000000000101000100011000000,
						cb148 = 32'b00000000000000000111110101110111,
						cb149 = 32'b00000000000001001010000010101000,
						cb150 = 32'b10000000000000010001111000000010,
						cb151 = 32'b10000000000000110011110111100010,
						cb152 = 32'b00000000000000011100101010100011,
						cb153 = 32'b00000000000010000110101000111000,
						cb154 = 32'b00000000000000000010011111110000,
						cb155 = 32'b00000000000000000010111011101111,
						cb156 = 32'b00000000000000001000100001001110,
						cb157 = 32'b00000000000000110010011110010000,
						cb158 = 32'b10000000000000001100001110110101,
						cb159 = 32'b00000000000100101000001110010101,
						cb160 = 32'b00000000000000001111001111010000,
						cb161 = 32'b00000000000010111100010101110011,
						cb162 = 32'b10000000000000000101010100100011,
						cb163 = 32'b00000000000000000101100011010100,
						cb164 = 32'b00000000000000000011001111000001,
						cb165 = 32'b00000000000011101011011110000000,
						cb166 = 32'b10000000000000100010000100010101,
						cb167 = 32'b10000000000011111000111100011010,
						cb168 = 32'b00000000000000010101101010000100,
						cb169 = 32'b10000000000000011110110101000010,
						cb170 = 32'b10000000000000000000001011001110,
						cb171 = 32'b10000000000100000101011000011110,
						cb172 = 32'b00000000000000000110011000101000,
						cb173 = 32'b10000000000000101100101001100010,
						cb174 = 32'b00000000000000001100000000101011,
						cb175 = 32'b00000000000111110010010111110110,
						cb176 = 32'b00000000000000001010011111011110,
						cb177 = 32'b00000000000110000111101101011101,
						cb178 = 32'b10000000000000000111010000000101,
						cb179 = 32'b10000000000000001011110001100010,
						cb180 = 32'b00000000000000000100100101110010,
						cb181 = 32'b00000000000001101000101111110100,
						cb182 = 32'b10000000000000001011011100110110,
						cb183 = 32'b10000000000011000101101110011000,
						cb184 = 32'b00000000000000011000110001101001,
						cb185 = 32'b00000000000000111101111101000110,
						cb186 = 32'b00000000000000000100010110011001,
						cb187 = 32'b00000000000000001100110101100110,
						cb188 = 32'b00000000000000001000000010000111,
						cb189 = 32'b10000000000001001101101011010111,
						cb190 = 32'b10000000000000000111111100111101,
						cb191 = 32'b00000000000100011100001100001011,
						cb192 = 32'b00000000000000010011000011101111,
						cb193 = 32'b00000000000011011111010001010011,
						cb194 = 32'b00000000000000000000010000000000,
						cb195 = 32'b00000000000000010101010011100001,
						cb196 = 32'b00000000000000000101011110000100,
						cb197 = 32'b00000000000010001110111101110100,
						cb198 = 32'b10000000000000100101000011100110,
						cb199 = 32'b10000000000001010110010100100010,
						cb200 = 32'b00000000000000001100001000110100,
						cb201 = 32'b00000000000000011111011011101001,
						cb202 = 32'b00000000000000000011110111000111,
						cb203 = 32'b10000000000000110011110011011001,
						cb204 = 32'b00000000000000000100010001100100,
						cb205 = 32'b10000000000010110011110000000001,
						cb206 = 32'b10000000000000000100010111101011,
						cb207 = 32'b00000000001000001001111111110010,
						cb208 = 32'b00000000000000011100000011100110,
						cb209 = 32'b00000000001010000110111010010111,
						cb210 = 32'b10000000000000001100100010110100,
						cb211 = 32'b00000000000000110000101110110110,
						cb212 = 32'b00000000000000001011010010111011,
						cb213 = 32'b00000000000001011010100101000011,
						cb214 = 32'b10000000000000010110001011101011,
						cb215 = 32'b00000000000000010101101010000010,
						cb216 = 32'b00000000000000100110000001011111,
						cb217 = 32'b00000000000000011010110011000010,
						cb218 = 32'b00000000000000000011111000110011,
						cb219 = 32'b00000000000001001011101101110000,
						cb220 = 32'b00000000000000000111110111000001,
						cb221 = 32'b00000000000000000101101010100011,
						cb222 = 32'b10000000000000011001101101010100,
						cb223 = 32'b00000000000010001010100010110000,
						cb224 = 32'b00000000000000010010101011000111,
						cb225 = 32'b00000000000001011111110010110010,
						cb226 = 32'b10000000000000000010001100111001,
						cb227 = 32'b10000000000011000000101010101100,
						cb228 = 32'b10000000000000000100000001011010,
						cb229 = 32'b00000000000010100110010110101110,
						cb230 = 32'b10000000000000010110111001110111,
						cb231 = 32'b10000000000010001110011101110011,
						cb232 = 32'b00000000000000001111110011111111,
						cb233 = 32'b10000000000011010011010110000001,
						cb234 = 32'b00000000000000000100001011110000,
						cb235 = 32'b10000000000001100101101011011111,
						cb236 = 32'b00000000000000000110010101011011,
						cb237 = 32'b10000000000000001011001111011000,
						cb238 = 32'b00000000000000000100100010100000,
						cb239 = 32'b00000000000110101110011001001100,
						cb240 = 32'b00000000000000000110101111000011,
						cb241 = 32'b00000000000011110111000100011001,
						cb242 = 32'b10000000000000000101101100010101,
						cb243 = 32'b10000000000011011011101001010001,
						cb244 = 32'b00000000000000001000011100000001,
						cb245 = 32'b00000000000011000110011000000100,
						cb246 = 32'b10000000000000010010101101101000,
						cb247 = 32'b10000000000011111111111110011101,
						cb248 = 32'b00000000000000011110100000011100,
						cb249 = 32'b10000000000001011101000011101000,
						cb250 = 32'b00000000000000000101101010111111,
						cb251 = 32'b00000000000000111101101000000000,
						cb252 = 32'b00000000000000001101001101100101,
						cb253 = 32'b10000000000001000010100110100010,
						cb254 = 32'b10000000000000000111110101111101,
						cb255 = 32'b00000000000011010000111010100100,
						cb256 = 32'b00000000000000100100000101111010,
						cb257 = 32'b00000000000011011000011011000010,
						cb258 = 32'b10000000000000000000000101000100,
						cb259 = 32'b10000000000000110011110010110100,
						cb260 = 32'b00000000000000000000011011010110,
						cb261 = 32'b00000000000001111101110111001111,
						cb262 = 32'b10000000000000011100111101110100,
						cb263 = 32'b10000000000000000111001110000000,
						cb264 = 32'b00000000000000010001010101110101,
						cb265 = 32'b10000000000000000010111100000001,
						cb266 = 32'b00000000000000000010001011000110,
						cb267 = 32'b10000000000000100100010000111110,
						cb268 = 32'b00000000000000000110000000110101,
						cb269 = 32'b10000000000001011000001100100010,
						cb270 = 32'b10000000000000011111011101101000,
						cb271 = 32'b00000000001001101010111011010010,
						cb272 = 32'b00000000000000011111101001011101,
						cb273 = 32'b00000000000110001001000011000100,
						cb274 = 32'b10000000000000001011010001100100,
						cb275 = 32'b00000000000001100101101111011010,
						cb276 = 32'b00000000000000000111101100010100,
						cb277 = 32'b00000000000001110000110100111111,
						cb278 = 32'b10000000000000001111100111110110,
						cb279 = 32'b10000000000000100110110000111000,
						cb280 = 32'b00000000000000101000000010001100,
						cb281 = 32'b00000000000001101100001001100100,
						cb282 = 32'b00000000000000000001010101100110,
						cb283 = 32'b00000000000000110100001001000000,
						cb284 = 32'b00000000000000001000101100101011,
						cb285 = 32'b00000000000000001110100011110110,
						cb286 = 32'b10000000000000010011101101100001,
						cb287 = 32'b00000000000101110001011101101100,
						cb288 = 32'b00000000000000001100100100010110,
						cb289 = 32'b00000000000011101100111010010111,
						cb290 = 32'b10000000000000000011011010101011,
						cb291 = 32'b00000000000000011011000000100000,
						cb292 = 32'b00000000000000000000000100110111,
						cb293 = 32'b00000000000100100010101111111011,
						cb294 = 32'b10000000000000011000110000010100,
						cb295 = 32'b10000000000100000001110111100110,
						cb296 = 32'b00000000000000011000000001000100,
						cb297 = 32'b10000000000000110100011111111000,
						cb298 = 32'b00000000000000000001010010000011,
						cb299 = 32'b10000000000001001010001001111101,
						cb300 = 32'b00000000000000000111101000000001,
						cb301 = 32'b10000000000000100010111001010001,
						cb302 = 32'b00000000000000000111000101000101,
						cb303 = 32'b00000000001010000100110111010010,
						cb304 = 32'b00000000000000010001001010100001,
						cb305 = 32'b00000000000110111001011110001101,
						cb306 = 32'b10000000000000001001100001000000,
						cb307 = 32'b10000000000001000010101010110100,
						cb308 = 32'b00000000000000000110110000100111,
						cb309 = 32'b00000000000001111001110110111000,
						cb310 = 32'b10000000000000001110110101110010,
						cb311 = 32'b10000000000001110100011000111111,
						cb312 = 32'b00000000000000011111110111011010,
						cb313 = 32'b00000000000000010100101111011110,
						cb314 = 32'b00000000000000000100101010010011,
						cb315 = 32'b00000000000000100110011000010110,
						cb316 = 32'b00000000000000001011100010011000,
						cb317 = 32'b10000000000000011111001101011011,
						cb318 = 32'b10000000000000001100110111100011,
						cb319 = 32'b00000000000110001110110111110011,
						cb320 = 32'b00000000000000011010010111111100,
						cb321 = 32'b00000000000100110001111010100100,
						cb322 = 32'b00000000000000000000111110010011,
						cb323 = 32'b10000000000000001001011100110100,
						cb324 = 32'b00000000000000000100010000011110,
						cb325 = 32'b00000000000010010001101001101110,
						cb326 = 32'b10000000000000011111010100011000,
						cb327 = 32'b10000000000000101110001001110101,
						cb328 = 32'b00000000000000010001110111101111,
						cb329 = 32'b00000000000000101010110000100010,
						cb330 = 32'b00000000000000000101101011000101,
						cb331 = 32'b10000000000000101011111110100000,
						cb332 = 32'b00000000000000000101010010101010,
						cb333 = 32'b10000000000011100010011111110110,
						cb334 = 32'b10000000000000001000011100100001,
						cb335 = 32'b00000000001001111001001101011010,
						cb336 = 32'b00000000000000001111110110111100,
						cb337 = 32'b00000000001010110011000111101011,
						cb338 = 32'b10000000000000001001011011110001,
						cb339 = 32'b00000000000000010100010011101001,
						cb340 = 32'b00000000000000001100100110010011,
						cb341 = 32'b00000000000010001011101100001111,
						cb342 = 32'b10000000000000010000001110001000,
						cb343 = 32'b00000000000000010000011001101010,
						cb344 = 32'b00000000000000101101001101001101,
						cb345 = 32'b00000000000000011110010100110111,
						cb346 = 32'b00000000000000000011110110101010,
						cb347 = 32'b00000000000000101011111011011101,
						cb348 = 32'b00000000000000000110110101011100,
						cb349 = 32'b00000000000000101000101101100001,
						cb350 = 32'b10000000000000011111001111111111,
						cb351 = 32'b00000000000011000011111001110110,
						cb352 = 32'b00000000000000010111001011011000,
						cb353 = 32'b00000000000011000000111110001010,
						cb354 = 32'b10000000000000000011010111100010,
						cb355 = 32'b10000000000000110110000100001010,
						cb356 = 32'b10000000000000000000111010000100,
						cb357 = 32'b00000000000010100011010000111001,
						cb358 = 32'b10000000000000011010011100000001,
						cb359 = 32'b10000000000001010001101001001101,
						cb360 = 32'b00000000000000010100101101110100,
						cb361 = 32'b10000000000011000100010101010011,
						cb362 = 32'b00000000000000000001110010010010,
						cb363 = 32'b10000000000010001010110100001001,
						cb364 = 32'b00000000000000000101001110011110,
						cb365 = 32'b10000000000000010010101011101001,
						cb366 = 32'b00000000000000000000010110010011,
						cb367 = 32'b00000000000111110010000000110100,
						cb368 = 32'b00000000000000000111010010010000,
						cb369 = 32'b00000000000101010111011111101001,
						cb370 = 32'b10000000000000000110000000011100,
						cb371 = 32'b10000000000000110101111100000111,
						cb372 = 32'b00000000000000000110010011000100,
						cb373 = 32'b00000000000010110100110101001111,
						cb374 = 32'b10000000000000001101100111111001,
						cb375 = 32'b10000000000100110110101000110110,
						cb376 = 32'b00000000000000100001101101100110,
						cb377 = 32'b10000000000000100011101010010110,
						cb378 = 32'b00000000000000000101111110001100,
						cb379 = 32'b00000000000000011110110010001111,
						cb380 = 32'b00000000000000001110001001101010,
						cb381 = 32'b10000000000000011011100001110111,
						cb382 = 32'b10000000000000001111100110100001,
						cb383 = 32'b00000000000010011101011100010010,
						cb384 = 32'b00000000000000100000000011011000,
						cb385 = 32'b00000000000100010110010100111000,
						cb386 = 32'b10000000000000000000100101110011,
						cb387 = 32'b10000000000000010001110010000010,
						cb388 = 32'b00000000000000000010011000000001,
						cb389 = 32'b00000000000001010110011001100100,
						cb390 = 32'b10000000000000011110101000010110,
						cb391 = 32'b00000000000001001100011000011001,
						cb392 = 32'b00000000000000010111001010101010,
						cb393 = 32'b00000000000000001000100110000000,
						cb394 = 32'b00000000000000000011000111101010,
						cb395 = 32'b10000000000000010000100111000110,
						cb396 = 32'b00000000000000000111111011101010,
						cb397 = 32'b10000000000010011111010001111100,
						cb398 = 32'b10000000000000010000111100011001,
						cb399 = 32'b00000000001000001111001001110101,
						cb400 = 32'b00000000000000100000001011011111,
						cb401 = 32'b00000000001000000111010001010011,
						cb402 = 32'b10000000000000000100111101000101,
						cb403 = 32'b00000000000001001011100000010111,
						cb404 = 32'b00000000000000000110111110100011,
						cb405 = 32'b00000000000001001010001010110001,
						cb406 = 32'b10000000000000010011110010110011,
						cb407 = 32'b10000000000000010100000100011000,
						cb408 = 32'b00000000000000100000010111010010,
						cb409 = 32'b00000000000010010110110110100111,
						cb410 = 32'b00000000000000000011000010111010,
						cb411 = 32'b00000000000000010111010111110101,
						cb412 = 32'b00000000000000000111101010100000,
						cb413 = 32'b00000000000000100111110000011011,
						cb414 = 32'b10000000000000010001010000010111,
						cb415 = 32'b00000000000100000011100011000001,
						cb416 = 32'b00000000000000010011010100100111,
						cb417 = 32'b00000000000010011010011101111010,
						cb418 = 32'b10000000000000000100001000010001,
						cb419 = 32'b10000000000000011010110000011111,
						cb420 = 32'b00000000000000000001001001100100,
						cb421 = 32'b00000000000011010110101001111110,
						cb422 = 32'b10000000000000011110000010010010,
						cb423 = 32'b10000000000100000001001001101110,
						cb424 = 32'b00000000000000010100101000100001,
						cb425 = 32'b10000000000001001101111100000101,
						cb426 = 32'b00000000000000000001000101010101,
						cb427 = 32'b10000000000011010111000101010100,
						cb428 = 32'b00000000000000000110111110000000,
						cb429 = 32'b10000000000001000010101001011110,
						cb430 = 32'b00000000000000000111011101010100,
						cb431 = 32'b00000000000111101001011011101001,
						cb432 = 32'b00000000000000001110011110100111,
						cb433 = 32'b00000000000101011001100100010110,
						cb434 = 32'b10000000000000001000010010110011,
						cb435 = 32'b10000000000000101000100000110100,
						cb436 = 32'b00000000000000000101011001011101,
						cb437 = 32'b00000000000001011010001100100011,
						cb438 = 32'b10000000000000001000111000010010,
						cb439 = 32'b10000000000100010110011010000111,
						cb440 = 32'b00000000000000011011000100011111,
						cb441 = 32'b00000000000000010010010101001111,
						cb442 = 32'b00000000000000000011101001011001,
						cb443 = 32'b00000000000000001110001110101000,
						cb444 = 32'b00000000000000001001011001011001,
						cb445 = 32'b10000000000001011011101011001111,
						cb446 = 32'b10000000000000000100001100011011,
						cb447 = 32'b00000000000100101010101010100110,
						cb448 = 32'b00000000000000010110010100100001,
						cb449 = 32'b00000000000100010000000010111110,
						cb450 = 32'b10000000000000000000010011100011,
						cb451 = 32'b00000000000001000100111011110001,
						cb452 = 32'b00000000000000000100110111100010,
						cb453 = 32'b00000000000011001010101101111110,
						cb454 = 32'b10000000000000100001001011110101,
						cb455 = 32'b10000000000001100111010111111001,
						cb456 = 32'b00000000000000001110101110101000,
						cb457 = 32'b00000000000000010011011010000100,
						cb458 = 32'b00000000000000000100100011110000,
						cb459 = 32'b10000000000000011100100100010100,
						cb460 = 32'b00000000000000000011010110110000,
						cb461 = 32'b10000000000100000000011000100100,
						cb462 = 32'b10000000000000001010001011010101,
						cb463 = 32'b00000000000111111001001110101001,
						cb464 = 32'b00000000000000010101100110010010,
						cb465 = 32'b00000000001000101010110101110000,
						cb466 = 32'b10000000000000001111100010111100,
						cb467 = 32'b00000000000001010100110100000101,
						cb468 = 32'b00000000000000001001011100011010,
						cb469 = 32'b00000000000001000111001100100000,
						cb470 = 32'b10000000000000011001000101011111,
						cb471 = 32'b00000000000000111001101000110110,
						cb472 = 32'b00000000000000100010010100111111,
						cb473 = 32'b00000000000001001000010001000011,
						cb474 = 32'b00000000000000000100101111001000,
						cb475 = 32'b00000000000001000001111011000011,
						cb476 = 32'b00000000000000000111000111111111,
						cb477 = 32'b00000000000000001101111001100111,
						cb478 = 32'b10000000000000010111000100100010,
						cb479 = 32'b00000000000011100010000011011110,
						cb480 = 32'b00000000000000010101101100010010,
						cb481 = 32'b00000000000001100000000111100100,
						cb482 = 32'b10000000000000000000001101000111,
						cb483 = 32'b10000000000001110111111100011111,
						cb484 = 32'b10000000000000000110111000010100,
						cb485 = 32'b00000000000010001000000000000111,
						cb486 = 32'b10000000000000010011010001100110,
						cb487 = 32'b10000000000001110001110011111110,
						cb488 = 32'b00000000000000010001100111011100,
						cb489 = 32'b10000000000001101101011000111001,
						cb490 = 32'b00000000000000000011001001001011,
						cb491 = 32'b10000000000001100011101111100111,
						cb492 = 32'b00000000000000000110111111001110,
						cb493 = 32'b10000000000000010010000100111001,
						cb494 = 32'b00000000000000000010010000011011,
						cb495 = 32'b00000000000101101101101011011010,
						cb496 = 32'b00000000000000000100101001110011,
						cb497 = 32'b00000000000100101100111110110111,
						cb498 = 32'b10000000000000001000011110001111,
						cb499 = 32'b10000000000001111011101110000101,
						cb500 = 32'b00000000000000001010001001100000,
						cb501 = 32'b00000000000010101100101000110000,
						cb502 = 32'b10000000000000010101010110110000,
						cb503 = 32'b10000000000101000101001101100111,
						cb504 = 32'b00000000000000011101000011001101,
						cb505 = 32'b10000000000000011110011100111111,
						cb506 = 32'b00000000000000000110010100010000,
						cb507 = 32'b00000000000000111100110000101110,
						cb508 = 32'b00000000000000001011101110010001,
						cb509 = 32'b10000000000010000010111100001110,
						cb510 = 32'b10000000000000001011110111000010,
						cb511 = 32'b00000000000010111100010010101111;



//------------------------------------------------------------------
//                 -- Module Instantiations --                  
//------------------------------------------------------------------
parameter [N-1:0] ge_coeff0 = 32'b00000000000000001100110011001100;
parameter [N-1:0] ge_coeff1 = 32'b00000000000000001110011001100110;

reg [N-1:0] w0,w1;
reg [N-1:0] x0,x1,in_lt1,in_lt2,add1,add2,add3,add4,mult1,mult2,mult3,
			mult4,in_logx1,in_logx2;
			
reg [N-1:0] e;

wire lt1;			
wire [N-1:0] out_add1,out_add2,out_mult1,out_mult2,out_logx1,out_logx2;

reg [N-1:0] err0,err1,fn_err0,fn_err1,fn_w0,fn_w1,cw_x0,cw_x1,cw_xq0,cw_xq1,in_x;
wire [N-1:0] nearest;
			
wire [N-1:0] cw_w0,cw_w1;
			
reg startcw,startfnw,startlog1,startlog2;
wire donecw,donefnw,donelog1,donelog2;

fplessthan #(Q,N) fplt1(in_lt1,in_lt2,lt1);
qadd #(Q,N) adder1(add1,add2,out_add1);
qadd #(Q,N) adder2(add3,add4,out_add2);

qmult #(Q,N) multiplier1(mult1,mult2,out_mult1);
qmult #(Q,N) multiplier2(mult3,mult4,out_mult2);

//log10 #(Q,N) calc_log10(in_logx,out_logx);

compute_weights_opt 		cw  		(startcw,clk,rst,cw_x0,cw_x1,cw_xq0,cw_xq1,cw_w0,cw_w1,donecw);
find_nearest_weighted 	fnw 		(startfnw,clk,rst,fn_err0,fn_err1,fn_w0,fn_w1,nearest,donefnw);
fp_log10 					fplog1		(startlog1,clk,rst,in_logx1,out_logx1,donelog1);
fp_log10 					fplog2		(startlog2,clk,rst,in_logx2,out_logx2,donelog2);

//------------------------------------------------------------------
//                 -- Begin Declarations & Coding --                  
//------------------------------------------------------------------

always@(posedge clk or negedge rst)     // Determine STATE
begin

	if (rst == 1'b0)
		STATE <= START;
	else
		STATE <= NEXT_STATE;

end


always@(*)                              // Determine NEXT_STATE
begin
	case(STATE)

	START:
	begin
		if(startewoe == 1'b1)
		begin
			NEXT_STATE = CHECK_E;
		end
		else
		begin
			NEXT_STATE = START;
		end
	end

	CHECK_E:
	begin
		NEXT_STATE = SET_E;
	end

	SET_E:
	begin
		NEXT_STATE = PRECALC1_X0;
	end

	PRECALC1_X0:
	begin
		NEXT_STATE = PRECALC2_X0;
	end

	PRECALC2_X0:
	begin
		if(donelog1)
		begin
			NEXT_STATE = PRE_CALC3_X0;
		end
		else
		begin
			NEXT_STATE = PRECALC2_X0;
		end
	end

	PRE_CALC3_X0:
	begin
		NEXT_STATE = CALC_X0;
	end

	CALC_X0:
	begin
		if(donelog2)
		begin
			NEXT_STATE = PRECALC_X1;
		end
		else
		begin
			NEXT_STATE = CALC_X0;
		end
	end

	PRECALC_X1:
	begin
		NEXT_STATE = CALC_X1;
	end

	CALC_X1:
	begin
		NEXT_STATE = SET_CW;
	end

	SET_CW:
	begin
		if(donecw)
		begin
			NEXT_STATE = CALC_CW;
		end
		else
		begin
			NEXT_STATE = SET_CW;
		end
	end

	CALC_CW:
	begin
		NEXT_STATE = PRECALC1_ERR;
	end

	PRECALC1_ERR:
	begin
		NEXT_STATE = PRECALC2_ERR;
	end

	PRECALC2_ERR:
	begin
		NEXT_STATE = CALC_ERR;
	end

	CALC_ERR:
	begin
		NEXT_STATE = SET_FNW;
	end

	SET_FNW:
	begin
		if(donefnw)
		begin
			NEXT_STATE = CALC_FNW;
		end
		else
		begin
			NEXT_STATE = SET_FNW;
		end
	end

	CALC_FNW:
	begin
		NEXT_STATE = XQ0_MULT;
	end
	
	XQ0_MULT:
	begin
		NEXT_STATE = XQ0_ADD;
	end
	
	XQ0_ADD:
	begin
		NEXT_STATE = SET_XQ0;
	end
	
	SET_XQ0:
	begin
		NEXT_STATE = DONE;
	end

	DONE:
	begin
		NEXT_STATE = START;
	end

	endcase
end


always@(posedge clk or negedge rst)     // Determine outputs
begin

	if (rst == 1'b0)
	begin
		e <= 32'b0;
		doneewoe <= 1'b0;

	end

	else
	begin
		case(STATE)

		START:
		begin
			startfnw <= 1'b0;
			startcw <= 1'b0;
			startlog1 <= 1'b0;
			startlog2 <= 1'b0;
			doneewoe <= 1'b0;
		end

		CHECK_E:
		begin
			in_lt1 <= in_e;
			in_lt2 <= 32'b0;
		end

		SET_E:
		begin
			if(lt1)
			begin
				e <= 32'b0;
			end
			else
			begin
				e <= in_e;
			end
		end

		PRECALC1_X0:
		begin
			mult1 <= model_wo;
			mult2 <= 32'b00000000000110010111011011111100;
			
			//check_e <= e;
			add1 <= e;
			add2 <= 32'b00000000000000000000000000000110;
		end

		PRECALC2_X0:
		begin
			//check_mult <= out_mult1;
			in_logx1 <= out_mult1;
			startlog1 <= 1'b1;
		end

		PRE_CALC3_X0:
		begin
			
			mult1 <= out_logx1;
			mult2 <= 32'b00000000000000110101001001101001;
			startlog1 <= 1'b0;
		end

		CALC_X0:
		begin
			x0 <= out_mult1;
			
			in_logx2 <= out_add1;
			//check_add1 <= out_add1;
			startlog2 <= 1'b1;
		end


		PRECALC_X1:
		begin
			mult1 <= 32'b00000000000010100000000000000000;
			mult2 <= out_logx2;
			//check_logx <= out_logx2;
			
			
			startlog2 <= 1'b0;
		end

		CALC_X1:
		begin
			x1 <= out_mult1;
			startcw <= 1'b1;
		end

		SET_CW:
		begin
			//check_x0 <= x0;
			//check_x1 <= x1;
			cw_x0  <= x0;
			cw_x1  <= x1;
			cw_xq0 <= xq0;
			cw_xq1 <= xq1;
			startcw <= 1'b0;
		end

		CALC_CW:
		begin
			w0 <= cw_w0;
			w1 <= cw_w1;
		end

		PRECALC1_ERR:
		begin
			mult1 <= ge_coeff0;
			mult2 <= xq0;
			mult3 <= ge_coeff1;
			mult4 <= xq1;
		end

		PRECALC2_ERR:
		begin
			add1 <= x0;
			add2 <= {(out_mult1[N-1] == 0)?1'b1:1'b0,out_mult1[N-2:0]};
			add3 <= x1;
			add4 <= {(out_mult2[N-1] == 0)?1'b1:1'b0,out_mult2[N-2:0]};
		end

		CALC_ERR:
		begin
			err0 <= out_add1;
			err1 <= out_add2;
			startfnw <= 1'b1;
		end

		SET_FNW:
		begin
			fn_err0 <= err0;
			fn_err1 <= err1;
			fn_w0   <= w0;
			fn_w1   <= w1;
			startfnw <= 1'b0;
		end

		CALC_FNW:
		begin
			out_n1 <= nearest;
		end
		
		XQ0_MULT:
		begin
			mult1 <= ge_coeff0;
			mult2 <= xq0;
			
			mult3 <= ge_coeff1;
			mult4 <= xq1;
		end
		
		XQ0_ADD:
		begin
			add1 <= out_mult1;
			add3 <= out_mult2;
			case( 2 * out_n1 )
				10'd0  :         add2 <= cb0;
				10'd2  :         add2 <= cb2;
				10'd4  :         add2 <= cb4;
				10'd6  :         add2 <= cb6;
				10'd8  :         add2 <= cb8;
				10'd10  :         add2 <= cb10;
				10'd12  :         add2 <= cb12;
				10'd14  :         add2 <= cb14;
				10'd16  :         add2 <= cb16;
				10'd18  :         add2 <= cb18;
				10'd20  :         add2 <= cb20;
				10'd22  :         add2 <= cb22;
				10'd24  :         add2 <= cb24;
				10'd26  :         add2 <= cb26;
				10'd28  :         add2 <= cb28;
				10'd30  :         add2 <= cb30;
				10'd32  :         add2 <= cb32;
				10'd34  :         add2 <= cb34;
				10'd36  :         add2 <= cb36;
				10'd38  :         add2 <= cb38;
				10'd40  :         add2 <= cb40;
				10'd42  :         add2 <= cb42;
				10'd44  :         add2 <= cb44;
				10'd46  :         add2 <= cb46;
				10'd48  :         add2 <= cb48;
				10'd50  :         add2 <= cb50;
				10'd52  :         add2 <= cb52;
				10'd54  :         add2 <= cb54;
				10'd56  :         add2 <= cb56;
				10'd58  :         add2 <= cb58;
				10'd60  :         add2 <= cb60;
				10'd62  :         add2 <= cb62;
				10'd64  :         add2 <= cb64;
				10'd66  :         add2 <= cb66;
				10'd68  :         add2 <= cb68;
				10'd70  :         add2 <= cb70;
				10'd72  :         add2 <= cb72;
				10'd74  :         add2 <= cb74;
				10'd76  :         add2 <= cb76;
				10'd78  :         add2 <= cb78;
				10'd80  :         add2 <= cb80;
				10'd82  :         add2 <= cb82;
				10'd84  :         add2 <= cb84;
				10'd86  :         add2 <= cb86;
				10'd88  :         add2 <= cb88;
				10'd90  :         add2 <= cb90;
				10'd92  :         add2 <= cb92;
				10'd94  :         add2 <= cb94;
				10'd96  :         add2 <= cb96;
				10'd98  :         add2 <= cb98;
				10'd100  :         add2 <= cb100;
				10'd102  :         add2 <= cb102;
				10'd104  :         add2 <= cb104;
				10'd106  :         add2 <= cb106;
				10'd108  :         add2 <= cb108;
				10'd110  :         add2 <= cb110;
				10'd112  :         add2 <= cb112;
				10'd114  :         add2 <= cb114;
				10'd116  :         add2 <= cb116;
				10'd118  :         add2 <= cb118;
				10'd120  :         add2 <= cb120;
				10'd122  :         add2 <= cb122;
				10'd124  :         add2 <= cb124;
				10'd126  :         add2 <= cb126;
				10'd128  :         add2 <= cb128;
				10'd130  :         add2 <= cb130;
				10'd132  :         add2 <= cb132;
				10'd134  :         add2 <= cb134;
				10'd136  :         add2 <= cb136;
				10'd138  :         add2 <= cb138;
				10'd140  :         add2 <= cb140;
				10'd142  :         add2 <= cb142;
				10'd144  :         add2 <= cb144;
				10'd146  :         add2 <= cb146;
				10'd148  :         add2 <= cb148;
				10'd150  :         add2 <= cb150;
				10'd152  :         add2 <= cb152;
				10'd154  :         add2 <= cb154;
				10'd156  :         add2 <= cb156;
				10'd158  :         add2 <= cb158;
				10'd160  :         add2 <= cb160;
				10'd162  :         add2 <= cb162;
				10'd164  :         add2 <= cb164;
				10'd166  :         add2 <= cb166;
				10'd168  :         add2 <= cb168;
				10'd170  :         add2 <= cb170;
				10'd172  :         add2 <= cb172;
				10'd174  :         add2 <= cb174;
				10'd176  :         add2 <= cb176;
				10'd178  :         add2 <= cb178;
				10'd180  :         add2 <= cb180;
				10'd182  :         add2 <= cb182;
				10'd184  :         add2 <= cb184;
				10'd186  :         add2 <= cb186;
				10'd188  :         add2 <= cb188;
				10'd190  :         add2 <= cb190;
				10'd192  :         add2 <= cb192;
				10'd194  :         add2 <= cb194;
				10'd196  :         add2 <= cb196;
				10'd198  :         add2 <= cb198;
				10'd200  :         add2 <= cb200;
				10'd202  :         add2 <= cb202;
				10'd204  :         add2 <= cb204;
				10'd206  :         add2 <= cb206;
				10'd208  :         add2 <= cb208;
				10'd210  :         add2 <= cb210;
				10'd212  :         add2 <= cb212;
				10'd214  :         add2 <= cb214;
				10'd216  :         add2 <= cb216;
				10'd218  :         add2 <= cb218;
				10'd220  :         add2 <= cb220;
				10'd222  :         add2 <= cb222;
				10'd224  :         add2 <= cb224;
				10'd226  :         add2 <= cb226;
				10'd228  :         add2 <= cb228;
				10'd230  :         add2 <= cb230;
				10'd232  :         add2 <= cb232;
				10'd234  :         add2 <= cb234;
				10'd236  :         add2 <= cb236;
				10'd238  :         add2 <= cb238;
				10'd240  :         add2 <= cb240;
				10'd242  :         add2 <= cb242;
				10'd244  :         add2 <= cb244;
				10'd246  :         add2 <= cb246;
				10'd248  :         add2 <= cb248;
				10'd250  :         add2 <= cb250;
				10'd252  :         add2 <= cb252;
				10'd254  :         add2 <= cb254;
				10'd256  :         add2 <= cb256;
				10'd258  :         add2 <= cb258;
				10'd260  :         add2 <= cb260;
				10'd262  :         add2 <= cb262;
				10'd264  :         add2 <= cb264;
				10'd266  :         add2 <= cb266;
				10'd268  :         add2 <= cb268;
				10'd270  :         add2 <= cb270;
				10'd272  :         add2 <= cb272;
				10'd274  :         add2 <= cb274;
				10'd276  :         add2 <= cb276;
				10'd278  :         add2 <= cb278;
				10'd280  :         add2 <= cb280;
				10'd282  :         add2 <= cb282;
				10'd284  :         add2 <= cb284;
				10'd286  :         add2 <= cb286;
				10'd288  :         add2 <= cb288;
				10'd290  :         add2 <= cb290;
				10'd292  :         add2 <= cb292;
				10'd294  :         add2 <= cb294;
				10'd296  :         add2 <= cb296;
				10'd298  :         add2 <= cb298;
				10'd300  :         add2 <= cb300;
				10'd302  :         add2 <= cb302;
				10'd304  :         add2 <= cb304;
				10'd306  :         add2 <= cb306;
				10'd308  :         add2 <= cb308;
				10'd310  :         add2 <= cb310;
				10'd312  :         add2 <= cb312;
				10'd314  :         add2 <= cb314;
				10'd316  :         add2 <= cb316;
				10'd318  :         add2 <= cb318;
				10'd320  :         add2 <= cb320;
				10'd322  :         add2 <= cb322;
				10'd324  :         add2 <= cb324;
				10'd326  :         add2 <= cb326;
				10'd328  :         add2 <= cb328;
				10'd330  :         add2 <= cb330;
				10'd332  :         add2 <= cb332;
				10'd334  :         add2 <= cb334;
				10'd336  :         add2 <= cb336;
				10'd338  :         add2 <= cb338;
				10'd340  :         add2 <= cb340;
				10'd342  :         add2 <= cb342;
				10'd344  :         add2 <= cb344;
				10'd346  :         add2 <= cb346;
				10'd348  :         add2 <= cb348;
				10'd350  :         add2 <= cb350;
				10'd352  :         add2 <= cb352;
				10'd354  :         add2 <= cb354;
				10'd356  :         add2 <= cb356;
				10'd358  :         add2 <= cb358;
				10'd360  :         add2 <= cb360;
				10'd362  :         add2 <= cb362;
				10'd364  :         add2 <= cb364;
				10'd366  :         add2 <= cb366;
				10'd368  :         add2 <= cb368;
				10'd370  :         add2 <= cb370;
				10'd372  :         add2 <= cb372;
				10'd374  :         add2 <= cb374;
				10'd376  :         add2 <= cb376;
				10'd378  :         add2 <= cb378;
				10'd380  :         add2 <= cb380;
				10'd382  :         add2 <= cb382;
				10'd384  :         add2 <= cb384;
				10'd386  :         add2 <= cb386;
				10'd388  :         add2 <= cb388;
				10'd390  :         add2 <= cb390;
				10'd392  :         add2 <= cb392;
				10'd394  :         add2 <= cb394;
				10'd396  :         add2 <= cb396;
				10'd398  :         add2 <= cb398;
				10'd400  :         add2 <= cb400;
				10'd402  :         add2 <= cb402;
				10'd404  :         add2 <= cb404;
				10'd406  :         add2 <= cb406;
				10'd408  :         add2 <= cb408;
				10'd410  :         add2 <= cb410;
				10'd412  :         add2 <= cb412;
				10'd414  :         add2 <= cb414;
				10'd416  :         add2 <= cb416;
				10'd418  :         add2 <= cb418;
				10'd420  :         add2 <= cb420;
				10'd422  :         add2 <= cb422;
				10'd424  :         add2 <= cb424;
				10'd426  :         add2 <= cb426;
				10'd428  :         add2 <= cb428;
				10'd430  :         add2 <= cb430;
				10'd432  :         add2 <= cb432;
				10'd434  :         add2 <= cb434;
				10'd436  :         add2 <= cb436;
				10'd438  :         add2 <= cb438;
				10'd440  :         add2 <= cb440;
				10'd442  :         add2 <= cb442;
				10'd444  :         add2 <= cb444;
				10'd446  :         add2 <= cb446;
				10'd448  :         add2 <= cb448;
				10'd450  :         add2 <= cb450;
				10'd452  :         add2 <= cb452;
				10'd454  :         add2 <= cb454;
				10'd456  :         add2 <= cb456;
				10'd458  :         add2 <= cb458;
				10'd460  :         add2 <= cb460;
				10'd462  :         add2 <= cb462;
				10'd464  :         add2 <= cb464;
				10'd466  :         add2 <= cb466;
				10'd468  :         add2 <= cb468;
				10'd470  :         add2 <= cb470;
				10'd472  :         add2 <= cb472;
				10'd474  :         add2 <= cb474;
				10'd476  :         add2 <= cb476;
				10'd478  :         add2 <= cb478;
				10'd480  :         add2 <= cb480;
				10'd482  :         add2 <= cb482;
				10'd484  :         add2 <= cb484;
				10'd486  :         add2 <= cb486;
				10'd488  :         add2 <= cb488;
				10'd490  :         add2 <= cb490;
				10'd492  :         add2 <= cb492;
				10'd494  :         add2 <= cb494;
				10'd496  :         add2 <= cb496;
				10'd498  :         add2 <= cb498;
				10'd500  :         add2 <= cb500;
				10'd502  :         add2 <= cb502;
				10'd504  :         add2 <= cb504;
				10'd506  :         add2 <= cb506;
				10'd508  :         add2 <= cb508;
				10'd510  :         add2 <= cb510;

			endcase
			
			case( (2 * out_n1) + 1 )
				10'd1  :         add4 <= cb1;
				10'd3  :         add4 <= cb3;
				10'd5  :         add4 <= cb5;
				10'd7  :         add4 <= cb7;
				10'd9  :         add4 <= cb9;
				10'd11  :         add4 <= cb11;
				10'd13  :         add4 <= cb13;
				10'd15  :         add4 <= cb15;
				10'd17  :         add4 <= cb17;
				10'd19  :         add4 <= cb19;
				10'd21  :         add4 <= cb21;
				10'd23  :         add4 <= cb23;
				10'd25  :         add4 <= cb25;
				10'd27  :         add4 <= cb27;
				10'd29  :         add4 <= cb29;
				10'd31  :         add4 <= cb31;
				10'd33  :         add4 <= cb33;
				10'd35  :         add4 <= cb35;
				10'd37  :         add4 <= cb37;
				10'd39  :         add4 <= cb39;
				10'd41  :         add4 <= cb41;
				10'd43  :         add4 <= cb43;
				10'd45  :         add4 <= cb45;
				10'd47  :         add4 <= cb47;
				10'd49  :         add4 <= cb49;
				10'd51  :         add4 <= cb51;
				10'd53  :         add4 <= cb53;
				10'd55  :         add4 <= cb55;
				10'd57  :         add4 <= cb57;
				10'd59  :         add4 <= cb59;
				10'd61  :         add4 <= cb61;
				10'd63  :         add4 <= cb63;
				10'd65  :         add4 <= cb65;
				10'd67  :         add4 <= cb67;
				10'd69  :         add4 <= cb69;
				10'd71  :         add4 <= cb71;
				10'd73  :         add4 <= cb73;
				10'd75  :         add4 <= cb75;
				10'd77  :         add4 <= cb77;
				10'd79  :         add4 <= cb79;
				10'd81  :         add4 <= cb81;
				10'd83  :         add4 <= cb83;
				10'd85  :         add4 <= cb85;
				10'd87  :         add4 <= cb87;
				10'd89  :         add4 <= cb89;
				10'd91  :         add4 <= cb91;
				10'd93  :         add4 <= cb93;
				10'd95  :         add4 <= cb95;
				10'd97  :         add4 <= cb97;
				10'd99  :         add4 <= cb99;
				10'd101  :         add4 <= cb101;
				10'd103  :         add4 <= cb103;
				10'd105  :         add4 <= cb105;
				10'd107  :         add4 <= cb107;
				10'd109  :         add4 <= cb109;
				10'd111  :         add4 <= cb111;
				10'd113  :         add4 <= cb113;
				10'd115  :         add4 <= cb115;
				10'd117  :         add4 <= cb117;
				10'd119  :         add4 <= cb119;
				10'd121  :         add4 <= cb121;
				10'd123  :         add4 <= cb123;
				10'd125  :         add4 <= cb125;
				10'd127  :         add4 <= cb127;
				10'd129  :         add4 <= cb129;
				10'd131  :         add4 <= cb131;
				10'd133  :         add4 <= cb133;
				10'd135  :         add4 <= cb135;
				10'd137  :         add4 <= cb137;
				10'd139  :         add4 <= cb139;
				10'd141  :         add4 <= cb141;
				10'd143  :         add4 <= cb143;
				10'd145  :         add4 <= cb145;
				10'd147  :         add4 <= cb147;
				10'd149  :         add4 <= cb149;
				10'd151  :         add4 <= cb151;
				10'd153  :         add4 <= cb153;
				10'd155  :         add4 <= cb155;
				10'd157  :         add4 <= cb157;
				10'd159  :         add4 <= cb159;
				10'd161  :         add4 <= cb161;
				10'd163  :         add4 <= cb163;
				10'd165  :         add4 <= cb165;
				10'd167  :         add4 <= cb167;
				10'd169  :         add4 <= cb169;
				10'd171  :         add4 <= cb171;
				10'd173  :         add4 <= cb173;
				10'd175  :         add4 <= cb175;
				10'd177  :         add4 <= cb177;
				10'd179  :         add4 <= cb179;
				10'd181  :         add4 <= cb181;
				10'd183  :         add4 <= cb183;
				10'd185  :         add4 <= cb185;
				10'd187  :         add4 <= cb187;
				10'd189  :         add4 <= cb189;
				10'd191  :         add4 <= cb191;
				10'd193  :         add4 <= cb193;
				10'd195  :         add4 <= cb195;
				10'd197  :         add4 <= cb197;
				10'd199  :         add4 <= cb199;
				10'd201  :         add4 <= cb201;
				10'd203  :         add4 <= cb203;
				10'd205  :         add4 <= cb205;
				10'd207  :         add4 <= cb207;
				10'd209  :         add4 <= cb209;
				10'd211  :         add4 <= cb211;
				10'd213  :         add4 <= cb213;
				10'd215  :         add4 <= cb215;
				10'd217  :         add4 <= cb217;
				10'd219  :         add4 <= cb219;
				10'd221  :         add4 <= cb221;
				10'd223  :         add4 <= cb223;
				10'd225  :         add4 <= cb225;
				10'd227  :         add4 <= cb227;
				10'd229  :         add4 <= cb229;
				10'd231  :         add4 <= cb231;
				10'd233  :         add4 <= cb233;
				10'd235  :         add4 <= cb235;
				10'd237  :         add4 <= cb237;
				10'd239  :         add4 <= cb239;
				10'd241  :         add4 <= cb241;
				10'd243  :         add4 <= cb243;
				10'd245  :         add4 <= cb245;
				10'd247  :         add4 <= cb247;
				10'd249  :         add4 <= cb249;
				10'd251  :         add4 <= cb251;
				10'd253  :         add4 <= cb253;
				10'd255  :         add4 <= cb255;
				10'd257  :         add4 <= cb257;
				10'd259  :         add4 <= cb259;
				10'd261  :         add4 <= cb261;
				10'd263  :         add4 <= cb263;
				10'd265  :         add4 <= cb265;
				10'd267  :         add4 <= cb267;
				10'd269  :         add4 <= cb269;
				10'd271  :         add4 <= cb271;
				10'd273  :         add4 <= cb273;
				10'd275  :         add4 <= cb275;
				10'd277  :         add4 <= cb277;
				10'd279  :         add4 <= cb279;
				10'd281  :         add4 <= cb281;
				10'd283  :         add4 <= cb283;
				10'd285  :         add4 <= cb285;
				10'd287  :         add4 <= cb287;
				10'd289  :         add4 <= cb289;
				10'd291  :         add4 <= cb291;
				10'd293  :         add4 <= cb293;
				10'd295  :         add4 <= cb295;
				10'd297  :         add4 <= cb297;
				10'd299  :         add4 <= cb299;
				10'd301  :         add4 <= cb301;
				10'd303  :         add4 <= cb303;
				10'd305  :         add4 <= cb305;
				10'd307  :         add4 <= cb307;
				10'd309  :         add4 <= cb309;
				10'd311  :         add4 <= cb311;
				10'd313  :         add4 <= cb313;
				10'd315  :         add4 <= cb315;
				10'd317  :         add4 <= cb317;
				10'd319  :         add4 <= cb319;
				10'd321  :         add4 <= cb321;
				10'd323  :         add4 <= cb323;
				10'd325  :         add4 <= cb325;
				10'd327  :         add4 <= cb327;
				10'd329  :         add4 <= cb329;
				10'd331  :         add4 <= cb331;
				10'd333  :         add4 <= cb333;
				10'd335  :         add4 <= cb335;
				10'd337  :         add4 <= cb337;
				10'd339  :         add4 <= cb339;
				10'd341  :         add4 <= cb341;
				10'd343  :         add4 <= cb343;
				10'd345  :         add4 <= cb345;
				10'd347  :         add4 <= cb347;
				10'd349  :         add4 <= cb349;
				10'd351  :         add4 <= cb351;
				10'd353  :         add4 <= cb353;
				10'd355  :         add4 <= cb355;
				10'd357  :         add4 <= cb357;
				10'd359  :         add4 <= cb359;
				10'd361  :         add4 <= cb361;
				10'd363  :         add4 <= cb363;
				10'd365  :         add4 <= cb365;
				10'd367  :         add4 <= cb367;
				10'd369  :         add4 <= cb369;
				10'd371  :         add4 <= cb371;
				10'd373  :         add4 <= cb373;
				10'd375  :         add4 <= cb375;
				10'd377  :         add4 <= cb377;
				10'd379  :         add4 <= cb379;
				10'd381  :         add4 <= cb381;
				10'd383  :         add4 <= cb383;
				10'd385  :         add4 <= cb385;
				10'd387  :         add4 <= cb387;
				10'd389  :         add4 <= cb389;
				10'd391  :         add4 <= cb391;
				10'd393  :         add4 <= cb393;
				10'd395  :         add4 <= cb395;
				10'd397  :         add4 <= cb397;
				10'd399  :         add4 <= cb399;
				10'd401  :         add4 <= cb401;
				10'd403  :         add4 <= cb403;
				10'd405  :         add4 <= cb405;
				10'd407  :         add4 <= cb407;
				10'd409  :         add4 <= cb409;
				10'd411  :         add4 <= cb411;
				10'd413  :         add4 <= cb413;
				10'd415  :         add4 <= cb415;
				10'd417  :         add4 <= cb417;
				10'd419  :         add4 <= cb419;
				10'd421  :         add4 <= cb421;
				10'd423  :         add4 <= cb423;
				10'd425  :         add4 <= cb425;
				10'd427  :         add4 <= cb427;
				10'd429  :         add4 <= cb429;
				10'd431  :         add4 <= cb431;
				10'd433  :         add4 <= cb433;
				10'd435  :         add4 <= cb435;
				10'd437  :         add4 <= cb437;
				10'd439  :         add4 <= cb439;
				10'd441  :         add4 <= cb441;
				10'd443  :         add4 <= cb443;
				10'd445  :         add4 <= cb445;
				10'd447  :         add4 <= cb447;
				10'd449  :         add4 <= cb449;
				10'd451  :         add4 <= cb451;
				10'd453  :         add4 <= cb453;
				10'd455  :         add4 <= cb455;
				10'd457  :         add4 <= cb457;
				10'd459  :         add4 <= cb459;
				10'd461  :         add4 <= cb461;
				10'd463  :         add4 <= cb463;
				10'd465  :         add4 <= cb465;
				10'd467  :         add4 <= cb467;
				10'd469  :         add4 <= cb469;
				10'd471  :         add4 <= cb471;
				10'd473  :         add4 <= cb473;
				10'd475  :         add4 <= cb475;
				10'd477  :         add4 <= cb477;
				10'd479  :         add4 <= cb479;
				10'd481  :         add4 <= cb481;
				10'd483  :         add4 <= cb483;
				10'd485  :         add4 <= cb485;
				10'd487  :         add4 <= cb487;
				10'd489  :         add4 <= cb489;
				10'd491  :         add4 <= cb491;
				10'd493  :         add4 <= cb493;
				10'd495  :         add4 <= cb495;
				10'd497  :         add4 <= cb497;
				10'd499  :         add4 <= cb499;
				10'd501  :         add4 <= cb501;
				10'd503  :         add4 <= cb503;
				10'd505  :         add4 <= cb505;
				10'd507  :         add4 <= cb507;
				10'd509  :         add4 <= cb509;
				10'd511  :         add4 <= cb511;

			endcase
		end
		
		SET_XQ0:
		begin
			out_xq0 <= out_add1;
			out_xq1 <= out_add2;
		end
		
		
		

		DONE:
		begin
			doneewoe <= 1'b1;
		end

		endcase
	end

end


endmodule