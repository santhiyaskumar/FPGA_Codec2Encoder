/*
* Module         - ROM_speech_w[[
* Top module     - cbselect
* Project        - CODEC2_ENCODE_2400
* Developer      - Santhiya S
* Date           - Mon Feb 04 15:19:31 2019
*
* Description    -
* Inputs         -

*32 bits fixed point representation
   S - E  - M
   1 - 15 - 16
*/
module ROM_speech_w_48(addr,dataout);

	parameter N = 48;
	input [9:0] addr;
	output reg [N-1:0] dataout;

	reg [N-1:0] w[319:0];
	
	always@(*)
	begin

				w[0]  =  48'b000000000000000000000000000000000000000000000000;
				w[1]  =  48'b000000000000000000000000000000000000000000000000;
				w[2]  =  48'b000000000000000000000000000000000000000000000000;
				w[3]  =  48'b000000000000000000000000000000000000000000000000;
				w[4]  =  48'b000000000000000000000000000000000000000000000000;
				w[5]  =  48'b000000000000000000000000000000000000000000000000;
				w[6]  =  48'b000000000000000000000000000000000000000000000000;
				w[7]  =  48'b000000000000000000000000000000000000000000000000;
				w[8]  =  48'b000000000000000000000000000000000000000000000000;
				w[9]  =  48'b000000000000000000000000000000000000000000000000;
				w[10]  =  48'b000000000000000000000000000000000000000000000000;
				w[11]  =  48'b000000000000000000000000000000000000000000000000;
				w[12]  =  48'b000000000000000000000000000000000000000000000000;
				w[13]  =  48'b000000000000000000000000000000000000000000000000;
				w[14]  =  48'b000000000000000000000000000000000000000000000000;
				w[15]  =  48'b000000000000000000000000000000000000000000000000;
				w[16]  =  48'b000000000000000000000000000000000000000000000000;
				w[17]  =  48'b000000000000000000000000000000000000000000000000;
				w[18]  =  48'b000000000000000000000000000000000000000000000000;
				w[19]  =  48'b000000000000000000000000000000000000000000000000;
				w[20]  =  48'b000000000000000000000000000000000000000000000000;
				w[21]  =  48'b000000000000000000000000000000000000000000000000;
				w[22]  =  48'b000000000000000000000000000000000000100101000110;
				w[23]  =  48'b000000000000000000000000000000000010010100010110;
				w[24]  =  48'b000000000000000000000000000000000101001101101110;
				w[25]  =  48'b000000000000000000000000000000001001010001000111;
				w[26]  =  48'b000000000000000000000000000000001110011110011000;
				w[27]  =  48'b000000000000000000000000000000010100110101011000;
				w[28]  =  48'b000000000000000000000000000000011100010101110111;
				w[29]  =  48'b000000000000000000000000000000100100111111100111;
				w[30]  =  48'b000000000000000000000000000000101110110010010110;
				w[31]  =  48'b000000000000000000000000000000111001101101101111;
				w[32]  =  48'b000000000000000000000000000001000101110001011100;
				w[33]  =  48'b000000000000000000000000000001010010111101000010;
				w[34]  =  48'b000000000000000000000000000001100001010000000111;
				w[35]  =  48'b000000000000000000000000000001110000101010001100;
				w[36]  =  48'b000000000000000000000000000010000001001010110001;
				w[37]  =  48'b000000000000000000000000000010010010110001010100;
				w[38]  =  48'b000000000000000000000000000010100101011101010000;
				w[39]  =  48'b000000000000000000000000000010111001001101111110;
				w[40]  =  48'b000000000000000000000000000011001110000010110100;
				w[41]  =  48'b000000000000000000000000000011100011111011000111;
				w[42]  =  48'b000000000000000000000000000011111010110110001001;
				w[43]  =  48'b000000000000000000000000000100010010110011001011;
				w[44]  =  48'b000000000000000000000000000100101011110001011001;
				w[45]  =  48'b000000000000000000000000000101000101110000000000;
				w[46]  =  48'b000000000000000000000000000101100000101110001010;
				w[47]  =  48'b000000000000000000000000000101111100101010111101;
				w[48]  =  48'b000000000000000000000000000110011001100101100000;
				w[49]  =  48'b000000000000000000000000000110110111011100110111;
				w[50]  =  48'b000000000000000000000000000111010110010000000001;
				w[51]  =  48'b000000000000000000000000000111110101111110000000;
				w[52]  =  48'b000000000000000000000000001000010110100101110000;
				w[53]  =  48'b000000000000000000000000001000111000000110001110;
				w[54]  =  48'b000000000000000000000000001001011010011110010100;
				w[55]  =  48'b000000000000000000000000001001111101101100111001;
				w[56]  =  48'b000000000000000000000000001010100001110000110100;
				w[57]  =  48'b000000000000000000000000001011000110101000111000;
				w[58]  =  48'b000000000000000000000000001011101100010011111010;
				w[59]  =  48'b000000000000000000000000001100010010110000101010;
				w[60]  =  48'b000000000000000000000000001100111001111101111001;
				w[61]  =  48'b000000000000000000000000001101100001111010010010;
				w[62]  =  48'b000000000000000000000000001110001010100100100101;
				w[63]  =  48'b000000000000000000000000001110110011111011011011;
				w[64]  =  48'b000000000000000000000000001111011101111101011101;
				w[65]  =  48'b000000000000000000000000010000001000101001010100;
				w[66]  =  48'b000000000000000000000000010000110011111101100111;
				w[67]  =  48'b000000000000000000000000010001011111111000111010;
				w[68]  =  48'b000000000000000000000000010010001100011001110010;
				w[69]  =  48'b000000000000000000000000010010111001011110110010;
				w[70]  =  48'b000000000000000000000000010011100111000110011011;
				w[71]  =  48'b000000000000000000000000010100010101001111001110;
				w[72]  =  48'b000000000000000000000000010101000011110111101100;
				w[73]  =  48'b000000000000000000000000010101110010111110010000;
				w[74]  =  48'b000000000000000000000000010110100010100001011010;
				w[75]  =  48'b000000000000000000000000010111010010011111100110;
				w[76]  =  48'b000000000000000000000000011000000010110111001111;
				w[77]  =  48'b000000000000000000000000011000110011100110110001;
				w[78]  =  48'b000000000000000000000000011001100100101100100110;
				w[79]  =  48'b000000000000000000000000011010010110000111000110;
				w[80]  =  48'b000000000000000000000000011011000111110100101001;
				w[81]  =  48'b000000000000000000000000011011111001110011101001;
				w[82]  =  48'b000000000000000000000000011100101100000010011101;
				w[83]  =  48'b000000000000000000000000011101011110011111011011;
				w[84]  =  48'b000000000000000000000000011110010001001000111011;
				w[85]  =  48'b000000000000000000000000011111000011111101010010;
				w[86]  =  48'b000000000000000000000000011111110110111010110100;
				w[87]  =  48'b000000000000000000000000100000101001111111111001;
				w[88]  =  48'b000000000000000000000000100001011101001010110101;
				w[89]  =  48'b000000000000000000000000100010010000011001111110;
				w[90]  =  48'b000000000000000000000000100011000011101011101000;
				w[91]  =  48'b000000000000000000000000100011110110111110000110;
				w[92]  =  48'b000000000000000000000000100100101010001111110000;
				w[93]  =  48'b000000000000000000000000100101011101011110111000;
				w[94]  =  48'b000000000000000000000000100110010000101001110101;
				w[95]  =  48'b000000000000000000000000100111000011101110111001;
				w[96]  =  48'b000000000000000000000000100111110110101100011101;
				w[97]  =  48'b000000000000000000000000101000101001100000110011;
				w[98]  =  48'b000000000000000000000000101001011100001010010010;
				w[99]  =  48'b000000000000000000000000101010001110100111010001;
				w[100]  =  48'b000000000000000000000000101011000000110110000100;
				w[101]  =  48'b000000000000000000000000101011110010110101000100;
				w[102]  =  48'b000000000000000000000000101100100100100010101001;
				w[103]  =  48'b000000000000000000000000101101010101111101001000;
				w[104]  =  48'b000000000000000000000000101110000111000010111101;
				w[105]  =  48'b000000000000000000000000101110110111110010011110;
				w[106]  =  48'b000000000000000000000000101111101000001010000111;
				w[107]  =  48'b000000000000000000000000110000011000001000010011;
				w[108]  =  48'b000000000000000000000000110001000111101011011110;
				w[109]  =  48'b000000000000000000000000110001110110110010000010;
				w[110]  =  48'b000000000000000000000000110010100101011010011110;
				w[111]  =  48'b000000000000000000000000110011010011100011010011;
				w[112]  =  48'b000000000000000000000000110100000001001010111100;
				w[113]  =  48'b000000000000000000000000110100101110001111111100;
				w[114]  =  48'b000000000000000000000000110101011010110000110100;
				w[115]  =  48'b000000000000000000000000110110000110101100000111;
				w[116]  =  48'b000000000000000000000000110110110010000000011001;
				w[117]  =  48'b000000000000000000000000110111011100101100010000;
				w[118]  =  48'b000000000000000000000000111000000110101110010011;
				w[119]  =  48'b000000000000000000000000111000110000000101001000;
				w[120]  =  48'b000000000000000000000000111001011000101111011010;
				w[121]  =  48'b000000000000000000000000111010000000101011110100;
				w[122]  =  48'b000000000000000000000000111010100111111001000011;
				w[123]  =  48'b000000000000000000000000111011001110010101110101;
				w[124]  =  48'b000000000000000000000000111011110100000000110110;
				w[125]  =  48'b000000000000000000000000111100011000111000111011;
				w[126]  =  48'b000000000000000000000000111100111100111100110101;
				w[127]  =  48'b000000000000000000000000111101100000001011011010;
				w[128]  =  48'b000000000000000000000000111110000010100011011111;
				w[129]  =  48'b000000000000000000000000111110100100000011111110;
				w[130]  =  48'b000000000000000000000000111111000100101011101101;
				w[131]  =  48'b000000000000000000000000111111100100011001101100;
				w[132]  =  48'b000000000000000000000001000000000011001100110110;
				w[133]  =  48'b000000000000000000000001000000100001000100001100;
				w[134]  =  48'b000000000000000000000001000000111101111110110000;
				w[135]  =  48'b000000000000000000000001000001011001111011100100;
				w[136]  =  48'b000000000000000000000001000001110100111001101110;
				w[137]  =  48'b000000000000000000000001000010001110111000010110;
				w[138]  =  48'b000000000000000000000001000010100111110110100010;
				w[139]  =  48'b000000000000000000000001000010111111110011100100;
				w[140]  =  48'b000000000000000000000001000011010110101110101000;
				w[141]  =  48'b000000000000000000000001000011101100100110111010;
				w[142]  =  48'b000000000000000000000001000100000001011011110000;
				w[143]  =  48'b000000000000000000000001000100010101001100011110;
				w[144]  =  48'b000000000000000000000001000100100111111000011010;
				w[145]  =  48'b000000000000000000000001000100111001011110111100;
				w[146]  =  48'b000000000000000000000001000101001001111111100010;
				w[147]  =  48'b000000000000000000000001000101011001011001101000;
				w[148]  =  48'b000000000000000000000001000101100111101100101100;
				w[149]  =  48'b000000000000000000000001000101110100111000010010;
				w[150]  =  48'b000000000000000000000001000110000000111011111110;
				w[151]  =  48'b000000000000000000000001000110001011110111011000;
				w[152]  =  48'b000000000000000000000001000110010101101010000110;
				w[153]  =  48'b000000000000000000000001000110011110010011110110;
				w[154]  =  48'b000000000000000000000001000110100101110100010110;
				w[155]  =  48'b000000000000000000000001000110101100001011010110;
				w[156]  =  48'b000000000000000000000001000110110001011000100110;
				w[157]  =  48'b000000000000000000000001000110110101011011111110;
				w[158]  =  48'b000000000000000000000001000110111000010101010110;
				w[159]  =  48'b000000000000000000000001000110111010000100101000;
				w[160]  =  48'b000000000000000000000001000110111010101001101110;
				w[161]  =  48'b000000000000000000000001000110111010000100101000;
				w[162]  =  48'b000000000000000000000001000110111000010101011000;
				w[163]  =  48'b000000000000000000000001000110110101011011111110;
				w[164]  =  48'b000000000000000000000001000110110001011000100110;
				w[165]  =  48'b000000000000000000000001000110101100001011010110;
				w[166]  =  48'b000000000000000000000001000110100101110100010110;
				w[167]  =  48'b000000000000000000000001000110011110010011110110;
				w[168]  =  48'b000000000000000000000001000110010101101010000110;
				w[169]  =  48'b000000000000000000000001000110001011110111011000;
				w[170]  =  48'b000000000000000000000001000110000000111011111110;
				w[171]  =  48'b000000000000000000000001000101110100111000010010;
				w[172]  =  48'b000000000000000000000001000101100111101100101100;
				w[173]  =  48'b000000000000000000000001000101011001011001100110;
				w[174]  =  48'b000000000000000000000001000101001001111111100010;
				w[175]  =  48'b000000000000000000000001000100111001011110111100;
				w[176]  =  48'b000000000000000000000001000100100111111000011010;
				w[177]  =  48'b000000000000000000000001000100010101001100011110;
				w[178]  =  48'b000000000000000000000001000100000001011011110000;
				w[179]  =  48'b000000000000000000000001000011101100100110111010;
				w[180]  =  48'b000000000000000000000001000011010110101110101000;
				w[181]  =  48'b000000000000000000000001000010111111110011100100;
				w[182]  =  48'b000000000000000000000001000010100111110110100010;
				w[183]  =  48'b000000000000000000000001000010001110111000010100;
				w[184]  =  48'b000000000000000000000001000001110100111001101110;
				w[185]  =  48'b000000000000000000000001000001011001111011100100;
				w[186]  =  48'b000000000000000000000001000000111101111110110000;
				w[187]  =  48'b000000000000000000000001000000100001000100001100;
				w[188]  =  48'b000000000000000000000001000000000011001100111000;
				w[189]  =  48'b000000000000000000000000111111100100011001101100;
				w[190]  =  48'b000000000000000000000000111111000100101011101101;
				w[191]  =  48'b000000000000000000000000111110100100000011111110;
				w[192]  =  48'b000000000000000000000000111110000010100011100000;
				w[193]  =  48'b000000000000000000000000111101100000001011011010;
				w[194]  =  48'b000000000000000000000000111100111100111100110110;
				w[195]  =  48'b000000000000000000000000111100011000111000111001;
				w[196]  =  48'b000000000000000000000000111011110100000000110101;
				w[197]  =  48'b000000000000000000000000111011001110010101110010;
				w[198]  =  48'b000000000000000000000000111010100111111001000011;
				w[199]  =  48'b000000000000000000000000111010000000101011110111;
				w[200]  =  48'b000000000000000000000000111001011000101111011011;
				w[201]  =  48'b000000000000000000000000111000110000000101000110;
				w[202]  =  48'b000000000000000000000000111000000110101110010011;
				w[203]  =  48'b000000000000000000000000110111011100101100001111;
				w[204]  =  48'b000000000000000000000000110110110010000000011011;
				w[205]  =  48'b000000000000000000000000110110000110101100000110;
				w[206]  =  48'b000000000000000000000000110101011010110000110100;
				w[207]  =  48'b000000000000000000000000110100101110001111111011;
				w[208]  =  48'b000000000000000000000000110100000001001010111101;
				w[209]  =  48'b000000000000000000000000110011010011100011010010;
				w[210]  =  48'b000000000000000000000000110010100101011010100001;
				w[211]  =  48'b000000000000000000000000110001110110110010000010;
				w[212]  =  48'b000000000000000000000000110001000111101011100000;
				w[213]  =  48'b000000000000000000000000110000011000001000010100;
				w[214]  =  48'b000000000000000000000000101111101000001010000110;
				w[215]  =  48'b000000000000000000000000101110110111110010011110;
				w[216]  =  48'b000000000000000000000000101110000111000010111011;
				w[217]  =  48'b000000000000000000000000101101010101111101001001;
				w[218]  =  48'b000000000000000000000000101100100100100010101000;
				w[219]  =  48'b000000000000000000000000101011110010110101000110;
				w[220]  =  48'b000000000000000000000000101011000000110110000011;
				w[221]  =  48'b000000000000000000000000101010001110100111010010;
				w[222]  =  48'b000000000000000000000000101001011100001010010010;
				w[223]  =  48'b000000000000000000000000101000101001100000110101;
				w[224]  =  48'b000000000000000000000000100111110110101100011100;
				w[225]  =  48'b000000000000000000000000100111000011101110111000;
				w[226]  =  48'b000000000000000000000000100110010000101001110101;
				w[227]  =  48'b000000000000000000000000100101011101011110110111;
				w[228]  =  48'b000000000000000000000000100100101010001111110000;
				w[229]  =  48'b000000000000000000000000100011110110111110000101;
				w[230]  =  48'b000000000000000000000000100011000011101011101001;
				w[231]  =  48'b000000000000000000000000100010010000011001111101;
				w[232]  =  48'b000000000000000000000000100001011101001010110111;
				w[233]  =  48'b000000000000000000000000100000101001111111111001;
				w[234]  =  48'b000000000000000000000000011111110110111010110110;
				w[235]  =  48'b000000000000000000000000011111000011111101010001;
				w[236]  =  48'b000000000000000000000000011110010001001000111101;
				w[237]  =  48'b000000000000000000000000011101011110011111011100;
				w[238]  =  48'b000000000000000000000000011100101100000010011011;
				w[239]  =  48'b000000000000000000000000011011111001110011101010;
				w[240]  =  48'b000000000000000000000000011011000111110100101000;
				w[241]  =  48'b000000000000000000000000011010010110000111000110;
				w[242]  =  48'b000000000000000000000000011001100100101100100101;
				w[243]  =  48'b000000000000000000000000011000110011100110110011;
				w[244]  =  48'b000000000000000000000000011000000010110111001111;
				w[245]  =  48'b000000000000000000000000010111010010011111101000;
				w[246]  =  48'b000000000000000000000000010110100010100001011010;
				w[247]  =  48'b000000000000000000000000010101110010111110010010;
				w[248]  =  48'b000000000000000000000000010101000011110111101011;
				w[249]  =  48'b000000000000000000000000010100010101001111001100;
				w[250]  =  48'b000000000000000000000000010011100111000110011100;
				w[251]  =  48'b000000000000000000000000010010111001011110110000;
				w[252]  =  48'b000000000000000000000000010010001100011001110011;
				w[253]  =  48'b000000000000000000000000010001011111111000111001;
				w[254]  =  48'b000000000000000000000000010000110011111101101000;
				w[255]  =  48'b000000000000000000000000010000001000101001010011;
				w[256]  =  48'b000000000000000000000000001111011101111101011110;
				w[257]  =  48'b000000000000000000000000001110110011111011011010;
				w[258]  =  48'b000000000000000000000000001110001010100100100111;
				w[259]  =  48'b000000000000000000000000001101100001111010010010;
				w[260]  =  48'b000000000000000000000000001100111001111101110111;
				w[261]  =  48'b000000000000000000000000001100010010110000101010;
				w[262]  =  48'b000000000000000000000000001011101100010011111001;
				w[263]  =  48'b000000000000000000000000001011000110101000111000;
				w[264]  =  48'b000000000000000000000000001010100001110000110010;
				w[265]  =  48'b000000000000000000000000001001111101101100111001;
				w[266]  =  48'b000000000000000000000000001001011010011110010011;
				w[267]  =  48'b000000000000000000000000001000111000000110001111;
				w[268]  =  48'b000000000000000000000000001000010110100101110000;
				w[269]  =  48'b000000000000000000000000000111110101111110000001;
				w[270]  =  48'b000000000000000000000000000111010110010000000001;
				w[271]  =  48'b000000000000000000000000000110110111011100111000;
				w[272]  =  48'b000000000000000000000000000110011001100101100000;
				w[273]  =  48'b000000000000000000000000000101111100101010111100;
				w[274]  =  48'b000000000000000000000000000101100000101110001010;
				w[275]  =  48'b000000000000000000000000000101000101101111111111;
				w[276]  =  48'b000000000000000000000000000100101011110001011010;
				w[277]  =  48'b000000000000000000000000000100010010110011001010;
				w[278]  =  48'b000000000000000000000000000011111010110110001010;
				w[279]  =  48'b000000000000000000000000000011100011111011000111;
				w[280]  =  48'b000000000000000000000000000011001110000010110101;
				w[281]  =  48'b000000000000000000000000000010111001001101111110;
				w[282]  =  48'b000000000000000000000000000010100101011101010000;
				w[283]  =  48'b000000000000000000000000000010010010110001010100;
				w[284]  =  48'b000000000000000000000000000010000001001010110000;
				w[285]  =  48'b000000000000000000000000000001110000101010001100;
				w[286]  =  48'b000000000000000000000000000001100001010000000110;
				w[287]  =  48'b000000000000000000000000000001010010111101000010;
				w[288]  =  48'b000000000000000000000000000001000101110001011011;
				w[289]  =  48'b000000000000000000000000000000111001101101101111;
				w[290]  =  48'b000000000000000000000000000000101110110010010110;
				w[291]  =  48'b000000000000000000000000000000100100111111101000;
				w[292]  =  48'b000000000000000000000000000000011100010101110111;
				w[293]  =  48'b000000000000000000000000000000010100110101011000;
				w[294]  =  48'b000000000000000000000000000000001110011110011000;
				w[295]  =  48'b000000000000000000000000000000001001010001000111;
				w[296]  =  48'b000000000000000000000000000000000101001101101110;
				w[297]  =  48'b000000000000000000000000000000000010010100010110;
				w[298]  =  48'b000000000000000000000000000000000000100101000110;
				w[299]  =  48'b000000000000000000000000000000000000000000000000;
				w[300]  =  48'b000000000000000000000000000000000000000000000000;
				w[301]  =  48'b000000000000000000000000000000000000000000000000;
				w[302]  =  48'b000000000000000000000000000000000000000000000000;
				w[303]  =  48'b000000000000000000000000000000000000000000000000;
				w[304]  =  48'b000000000000000000000000000000000000000000000000;
				w[305]  =  48'b000000000000000000000000000000000000000000000000;
				w[306]  =  48'b000000000000000000000000000000000000000000000000;
				w[307]  =  48'b000000000000000000000000000000000000000000000000;
				w[308]  =  48'b000000000000000000000000000000000000000000000000;
				w[309]  =  48'b000000000000000000000000000000000000000000000000;
				w[310]  =  48'b000000000000000000000000000000000000000000000000;
				w[311]  =  48'b000000000000000000000000000000000000000000000000;
				w[312]  =  48'b000000000000000000000000000000000000000000000000;
				w[313]  =  48'b000000000000000000000000000000000000000000000000;
				w[314]  =  48'b000000000000000000000000000000000000000000000000;
				w[315]  =  48'b000000000000000000000000000000000000000000000000;
				w[316]  =  48'b000000000000000000000000000000000000000000000000;
				w[317]  =  48'b000000000000000000000000000000000000000000000000;
				w[318]  =  48'b000000000000000000000000000000000000000000000000;
				w[319]  =  48'b000000000000000000000000000000000000000000000000;
	
	
	
		dataout = w[addr];
	end
endmodule
