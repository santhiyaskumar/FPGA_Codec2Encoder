/*
* Module         - ROM_cb2
* Top module     - cbselect
* Project        - CODEC2_ENCODE_2400
* Developer      - Santhiya S
* Date           - Mon Feb 04 15:19:31 2019
*
* Description    -
* Inputs         -
*static const float codes2[] = {
		500,
		550,
		600,
		650,
		700,
		750,
		800,
		850,
		900,
		950,
		1000,
		1050,
		1100,
		1150,
		1200,
		1250
*};
*32 bits fixed point representation
   S - E  - M
   1 - 15 - 16
*/
module ROM_cb2(addr,dataout);

	parameter N = 32;
	input [3:0] addr;
	//input CS;
	output reg [N-1:0] dataout;

	reg [N-1:0] cb2[15:0];
	
	always@(*)
	begin
			cb2[0] = 32'b00000001111101000000000000000000;
			cb2[1] = 32'b00000010001001100000000000000000;
			cb2[2] = 32'b00000010010110000000000000000000;
			cb2[3] = 32'b00000010100010100000000000000000;
			cb2[4] = 32'b00000010101111000000000000000000;
			cb2[5] = 32'b00000010111011100000000000000000;
			cb2[6] = 32'b00000011001000000000000000000000;
			cb2[7] = 32'b00000011010100100000000000000000;
			cb2[8] = 32'b00000011100001000000000000000000;
			cb2[9] = 32'b00000011101101100000000000000000;
			cb2[10] = 32'b00000011111010000000000000000000;
			cb2[11] = 32'b00000100000110100000000000000000;
			cb2[12] = 32'b00000100010011000000000000000000;
			cb2[13] = 32'b00000100011111100000000000000000;
			cb2[14] = 32'b00000100101100000000000000000000;
			cb2[15] = 32'b00000100111000100000000000000000;
		
		dataout = cb2[addr];
	end
endmodule
