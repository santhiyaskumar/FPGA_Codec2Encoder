/*
* Module         - ROM_cb0
* Top module     - cbselect
* Project        - CODEC2_ENCODE_2400
* Developer      - Santhiya S
* Date           - Mon Feb 04 15:19:31 2019
*
* Description    -
* Inputs         -
*static const float codes0[] = {
  225,
  250,
  275,
  300,
  325,
  350,
  375,
  400,
  425,
  450,
  475,
  500,
  525,
  550,
  575,
  600
*};
*32 bits fixed point representation
   S - E  - M
   1 - 15 - 16
*/
module ROM_cb0(addr,dataout);

	parameter N = 32;
	input [3:0] addr;
	output reg [N-1:0] dataout;

	reg [N-1:0] cb0[15:0];
	
	always@(*)
	begin
		cb0[0] = 32'b00000000111000010000000000000000;
		cb0[1] = 32'b00000000111110100000000000000000;
		cb0[2] = 32'b00000001000100110000000000000000;
		cb0[3] = 32'b00000001001011000000000000000000;
		cb0[4] = 32'b00000001010001010000000000000000;
		cb0[5] = 32'b00000001010111100000000000000000;
		cb0[6] = 32'b00000001011101110000000000000000;
		cb0[7] = 32'b00000001100100000000000000000000;
		cb0[8] = 32'b00000001101010010000000000000000;
		cb0[9] = 32'b00000001110000100000000000000000;
		cb0[10] = 32'b00000001110110110000000000000000;
		cb0[11] = 32'b00000001111101000000000000000000;
		cb0[12] = 32'b00000010000011010000000000000000;
		cb0[13] = 32'b00000010001001100000000000000000;
		cb0[14] = 32'b00000010001111110000000000000000;
		cb0[15] = 32'b00000010010110000000000000000000;
		
		dataout = cb0[addr];
	end
endmodule
