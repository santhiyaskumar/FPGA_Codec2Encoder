/*
* Module         - ROM_cb0
* Top module     - cbselect
* Project        - CODEC2_ENCODE_2400
* Developer      - Santhiya S
* Date           - Mon Feb 04 15:19:31 2019
*
* Description    -
* Inputs         -

*32 bits fixed point representation
   S - E  - M
   1 - 15 - 16
*/
module ROM_nlp_w(addr,dataout);

	parameter N = 80;
	input [5:0] addr;
	output reg [N-1:0] dataout;

	reg [N-1:0] nlp_w[63:0];
	
	always@(*)
	begin
nlp_w[0] = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
nlp_w[1] = 80'b00000000000000000000000000000000000000000000000000000000000000000000000010100010;
nlp_w[2] = 80'b00000000000000000000000000000000000000000000000000000000000000000000001010001001;
nlp_w[3] = 80'b00000000000000000000000000000000000000000000000000000000000000000000010110101111;
nlp_w[4] = 80'b00000000000000000000000000000000000000000000000000000000000000000000101000001101;
nlp_w[5] = 80'b00000000000000000000000000000000000000000000000000000000000000000000111110010110;
nlp_w[6] = 80'b00000000000000000000000000000000000000000000000000000000000000000001011000111101;
nlp_w[7] = 80'b00000000000000000000000000000000000000000000000000000000000000000001110111110010;
nlp_w[8] = 80'b00000000000000000000000000000000000000000000000000000000000000000010011010100000;
nlp_w[9] = 80'b00000000000000000000000000000000000000000000000000000000000000000011000000110001;
nlp_w[10] = 80'b00000000000000000000000000000000000000000000000000000000000000000011101010001101;
nlp_w[11] = 80'b00000000000000000000000000000000000000000000000000000000000000000100010110011010;
nlp_w[12] = 80'b00000000000000000000000000000000000000000000000000000000000000000101000100111100;
nlp_w[13] = 80'b00000000000000000000000000000000000000000000000000000000000000000101110101010101;
nlp_w[14] = 80'b00000000000000000000000000000000000000000000000000000000000000000110100111000101;
nlp_w[15] = 80'b00000000000000000000000000000000000000000000000000000000000000000111011001101111;
nlp_w[16] = 80'b00000000000000000000000000000000000000000000000000000000000000001000001100110000;
nlp_w[17] = 80'b00000000000000000000000000000000000000000000000000000000000000001000111111101010;
nlp_w[18] = 80'b00000000000000000000000000000000000000000000000000000000000000001001110001111011;
nlp_w[19] = 80'b00000000000000000000000000000000000000000000000000000000000000001010100011000100;
nlp_w[20] = 80'b00000000000000000000000000000000000000000000000000000000000000001011010010100101;
nlp_w[21] = 80'b00000000000000000000000000000000000000000000000000000000000000001100000000000000;
nlp_w[22] = 80'b00000000000000000000000000000000000000000000000000000000000000001100101010111000;
nlp_w[23] = 80'b00000000000000000000000000000000000000000000000000000000000000001101010010110010;
nlp_w[24] = 80'b00000000000000000000000000000000000000000000000000000000000000001101110111010100;
nlp_w[25] = 80'b00000000000000000000000000000000000000000000000000000000000000001110011000001000;
nlp_w[26] = 80'b00000000000000000000000000000000000000000000000000000000000000001110110100111000;
nlp_w[27] = 80'b00000000000000000000000000000000000000000000000000000000000000001111001101010010;
nlp_w[28] = 80'b00000000000000000000000000000000000000000000000000000000000000001111100001000111;
nlp_w[29] = 80'b00000000000000000000000000000000000000000000000000000000000000001111110000001010;
nlp_w[30] = 80'b00000000000000000000000000000000000000000000000000000000000000001111111010010010;
nlp_w[31] = 80'b00000000000000000000000000000000000000000000000000000000000000001111111111010111;
nlp_w[32] = 80'b00000000000000000000000000000000000000000000000000000000000000001111111111010111;
nlp_w[33] = 80'b00000000000000000000000000000000000000000000000000000000000000001111111010010010;
nlp_w[34] = 80'b00000000000000000000000000000000000000000000000000000000000000001111110000001010;
nlp_w[35] = 80'b00000000000000000000000000000000000000000000000000000000000000001111100001000111;
nlp_w[36] = 80'b00000000000000000000000000000000000000000000000000000000000000001111001101010010;
nlp_w[37] = 80'b00000000000000000000000000000000000000000000000000000000000000001110110100111000;
nlp_w[38] = 80'b00000000000000000000000000000000000000000000000000000000000000001110011000001000;
nlp_w[39] = 80'b00000000000000000000000000000000000000000000000000000000000000001101110111010100;
nlp_w[40] = 80'b00000000000000000000000000000000000000000000000000000000000000001101010010110010;
nlp_w[41] = 80'b00000000000000000000000000000000000000000000000000000000000000001100101010111000;
nlp_w[42] = 80'b00000000000000000000000000000000000000000000000000000000000000001011111111111111;
nlp_w[43] = 80'b00000000000000000000000000000000000000000000000000000000000000001011010010100101;
nlp_w[44] = 80'b00000000000000000000000000000000000000000000000000000000000000001010100011000100;
nlp_w[45] = 80'b00000000000000000000000000000000000000000000000000000000000000001001110001111011;
nlp_w[46] = 80'b00000000000000000000000000000000000000000000000000000000000000001000111111101010;
nlp_w[47] = 80'b00000000000000000000000000000000000000000000000000000000000000001000001100110000;
nlp_w[48] = 80'b00000000000000000000000000000000000000000000000000000000000000000111011001101111;
nlp_w[49] = 80'b00000000000000000000000000000000000000000000000000000000000000000110100111000101;
nlp_w[50] = 80'b00000000000000000000000000000000000000000000000000000000000000000101110101010101;
nlp_w[51] = 80'b00000000000000000000000000000000000000000000000000000000000000000101000100111100;
nlp_w[52] = 80'b00000000000000000000000000000000000000000000000000000000000000000100010110011010;
nlp_w[53] = 80'b00000000000000000000000000000000000000000000000000000000000000000011101010001101;
nlp_w[54] = 80'b00000000000000000000000000000000000000000000000000000000000000000011000000110001;
nlp_w[55] = 80'b00000000000000000000000000000000000000000000000000000000000000000010011010100000;
nlp_w[56] = 80'b00000000000000000000000000000000000000000000000000000000000000000001110111110010;
nlp_w[57] = 80'b00000000000000000000000000000000000000000000000000000000000000000001011000111101;
nlp_w[58] = 80'b00000000000000000000000000000000000000000000000000000000000000000000111110010110;
nlp_w[59] = 80'b00000000000000000000000000000000000000000000000000000000000000000000101000001101;
nlp_w[60] = 80'b00000000000000000000000000000000000000000000000000000000000000000000010110101111;
nlp_w[61] = 80'b00000000000000000000000000000000000000000000000000000000000000000000001010001001;
nlp_w[62] = 80'b00000000000000000000000000000000000000000000000000000000000000000000000010100010;
nlp_w[63] = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
		
		dataout = nlp_w[addr];
	end
endmodule
