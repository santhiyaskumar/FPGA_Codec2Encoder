module parameter_test();
 
//   input clk;
//	output reg [7:0] out;  
//	
//	parameter [7:0] cb [0:7] = {8d'0,8d'1,8d'2,8d'3,8d'4,8d'5,8d'6,8d'7};
//	
//	reg [2:0] j = 3'b0;
//	
//	always@(posedge clk)
//	begin
//		if(j < 8) 
//		begin
//			j <= j+1;
//			out <= cb[j];
//		end
//		else
//		begin
//			j <= 0;
//			out <= 0;
//		end
//	end
//	
	


endmodule