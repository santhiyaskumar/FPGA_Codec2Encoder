/*
* Module 		- quantise
* Top module	- encode_lsps_scalar
* CODEC2_ENCODE_2400

Description: Compute the vector index
Inputs : m,k,cb[],vec[],w[],se

*32 bits fixed point representation

S - E	 - M
1 - 15 - 16

Simulation - Waveform16.vwf
*/

module quantise (clk,rst,startq,m,orderi,vec,besti,doneq);

//------------------------------------------------------------------
//                 -- Input/Output Declarations --                  
//------------------------------------------------------------------

	parameter N = 32;
	parameter Q = 16;
	
	input clk, rst;
	input startq;
	input [4:0] m;
	input [3:0] orderi;
	input [N-1:0] vec;
	
	output reg [4:0] besti;
	output reg doneq;
	reg [N-1:0] e;
	
	reg [N-1:0] beste;
	reg [N-1:0] cb0,cb1,cb2,cb3,cb4,cb5,cb6,cb7,cb8,cb9,cb10,cb11,cb12,cb13,cb14,cb15;
	reg [N-1:0] in_e,in_beste;
	reg [4:0] j;
	
	reg [N-1:0] in_e1,in_e2;
	reg [N-1:0] abs_e;
	wire [N-1:0] power_e;
	
	wire [N-1:0] out_e0,out_e1,out_e2,out_e3,out_e4,out_e5,out_e6,out_e7,out_e8,out_e9,out_e10,
					 out_e11,out_e12,out_e13,out_e14,out_e15;
	wire lt1;
	
	
	//reg [N-1:0] neg_vec = {(vec[N-1] == 0)?1'b1:1'b0,vec[N-2:0]};
	
// Cb values
parameter [N-1:0] cb0_0 = 32'b00000000111000010000000000000000,
						cb0_1 = 32'b00000000111110100000000000000000,
						cb0_2 = 32'b00000001000100110000000000000000,
						cb0_3 = 32'b00000001001011000000000000000000,
						cb0_4 = 32'b00000001010001010000000000000000,
						cb0_5 = 32'b00000001010111100000000000000000,
						cb0_6 = 32'b00000001011101110000000000000000,
						cb0_7 = 32'b00000001100100000000000000000000,
						cb0_8 = 32'b00000001101010010000000000000000,
						cb0_9 = 32'b00000001110000100000000000000000,
						cb0_10 = 32'b00000001110110110000000000000000,
						cb0_11 = 32'b00000001111101000000000000000000,
						cb0_12 = 32'b00000010000011010000000000000000,
						cb0_13 = 32'b00000010001001100000000000000000,
						cb0_14 = 32'b00000010001111110000000000000000,
						cb0_15 = 32'b00000010010110000000000000000000,
						
						cb1_0 = 32'b00000001010001010000000000000000,
						cb1_1 = 32'b00000001010111100000000000000000,
						cb1_2 = 32'b00000001011101110000000000000000,
						cb1_3 = 32'b00000001100100000000000000000000,
						cb1_4 = 32'b00000001101010010000000000000000,
						cb1_5 = 32'b00000001110000100000000000000000,
						cb1_6 = 32'b00000001110110110000000000000000,
						cb1_7 = 32'b00000001111101000000000000000000,
						cb1_8 = 32'b00000010000011010000000000000000,
						cb1_9 = 32'b00000010001001100000000000000000,
						cb1_10 = 32'b00000010001111110000000000000000,
						cb1_11 = 32'b00000010010110000000000000000000,
						cb1_12 = 32'b00000010011100010000000000000000,
						cb1_13 = 32'b00000010100010100000000000000000,
						cb1_14 = 32'b00000010101000110000000000000000,
						cb1_15 = 32'b00000010101111000000000000000000,
						
						cb2_0 = 32'b00000001111101000000000000000000,
						cb2_1 = 32'b00000010001001100000000000000000,
						cb2_2 = 32'b00000010010110000000000000000000,
						cb2_3 = 32'b00000010100010100000000000000000,
						cb2_4 = 32'b00000010101111000000000000000000,
						cb2_5 = 32'b00000010111011100000000000000000,
						cb2_6 = 32'b00000011001000000000000000000000,
						cb2_7 = 32'b00000011010100100000000000000000,
						cb2_8 = 32'b00000011100001000000000000000000,
						cb2_9 = 32'b00000011101101100000000000000000,
						cb2_10 = 32'b00000011111010000000000000000000,
						cb2_11 = 32'b00000100000110100000000000000000,
						cb2_12 = 32'b00000100010011000000000000000000,
						cb2_13 = 32'b00000100011111100000000000000000,
						cb2_14 = 32'b00000100101100000000000000000000,
						cb2_15 = 32'b00000100111000100000000000000000,
						
						cb3_0 = 32'b00000010101111000000000000000000,
						cb3_1 = 32'b00000011001000000000000000000000,
						cb3_2 = 32'b00000011100001000000000000000000,
						cb3_3 = 32'b00000011111010000000000000000000,
						cb3_4 = 32'b00000100010011000000000000000000,
						cb3_5 = 32'b00000100101100000000000000000000,
						cb3_6 = 32'b00000101000101000000000000000000,
						cb3_7 = 32'b00000101011110000000000000000000,
						cb3_8 = 32'b00000101110111000000000000000000,
						cb3_9 = 32'b00000110010000000000000000000000,
						cb3_10 = 32'b00000110101001000000000000000000,
						cb3_11 = 32'b00000111000010000000000000000000,
						cb3_12 = 32'b00000111011011000000000000000000,
						cb3_13 = 32'b00000111110100000000000000000000,
						cb3_14 = 32'b00001000001101000000000000000000,
						cb3_15 = 32'b00001000100110000000000000000000,
						
						cb4_0 = 32'b00000011101101100000000000000000,
						cb4_1 = 32'b00000100000110100000000000000000,
						cb4_2 = 32'b00000100011111100000000000000000,
						cb4_3 = 32'b00000100111000100000000000000000,
						cb4_4 = 32'b00000101010001100000000000000000,
						cb4_5 = 32'b00000101101010100000000000000000,
						cb4_6 = 32'b00000110000011100000000000000000,
						cb4_7 = 32'b00000110011100100000000000000000,
						cb4_8 = 32'b00000110110101100000000000000000,
						cb4_9 = 32'b00000111001110100000000000000000,
						cb4_10 = 32'b00000111100111100000000000000000,
						cb4_11 = 32'b00001000000000100000000000000000,
						cb4_12 = 32'b00001000011001100000000000000000,
						cb4_13 = 32'b00001000110010100000000000000000,
						cb4_14 = 32'b00001001001011100000000000000000,
						cb4_15 = 32'b00001001100100100000000000000000,
						
						cb5_0 = 32'b00000100010011000000000000000000,
						cb5_1 = 32'b00000100101100000000000000000000,
						cb5_2 = 32'b00000101000101000000000000000000,
						cb5_3 = 32'b00000101011110000000000000000000,
						cb5_4 = 32'b00000101110111000000000000000000,
						cb5_5 = 32'b00000110010000000000000000000000,
						cb5_6 = 32'b00000110101001000000000000000000,
						cb5_7 = 32'b00000111000010000000000000000000,
						cb5_8 = 32'b00000111011011000000000000000000,
						cb5_9 = 32'b00000111110100000000000000000000,
						cb5_10 = 32'b00001000001101000000000000000000,
						cb5_11 = 32'b00001000100110000000000000000000,
						cb5_12 = 32'b00001000111111000000000000000000,
						cb5_13 = 32'b00001001011000000000000000000000,
						cb5_14 = 32'b00001001110001000000000000000000,
						cb5_15 = 32'b00001010001010000000000000000000,
						
						cb6_0 = 32'b00000101110111000000000000000000,
						cb6_1 = 32'b00000110010000000000000000000000,
						cb6_2 = 32'b00000110101001000000000000000000,
						cb6_3 = 32'b00000111000010000000000000000000,
						cb6_4 = 32'b00000111011011000000000000000000,
						cb6_5 = 32'b00000111110100000000000000000000,
						cb6_6 = 32'b00001000001101000000000000000000,
						cb6_7 = 32'b00001000100110000000000000000000,
						cb6_8 = 32'b00001000111111000000000000000000,
						cb6_9 = 32'b00001001011000000000000000000000,
						cb6_10 = 32'b00001001110001000000000000000000,
						cb6_11 = 32'b00001010001010000000000000000000,
						cb6_12 = 32'b00001010100011000000000000000000,
						cb6_13 = 32'b00001010111100000000000000000000,
						cb6_14 = 32'b00001011010101000000000000000000,
						cb6_15 = 32'b00001011101110000000000000000000,
						
						cb7_0 = 32'b00001000111111000000000000000000,
						cb7_1 = 32'b00001001011000000000000000000000,
						cb7_2 = 32'b00001001110001000000000000000000,
						cb7_3 = 32'b00001010001010000000000000000000,
						cb7_4 = 32'b00001010100011000000000000000000,
						cb7_5 = 32'b00001010111100000000000000000000,
						cb7_6 = 32'b00001011010101000000000000000000,
						cb7_7 = 32'b00001011101110000000000000000000,
						
						cb8_0 = 32'b00001001110001000000000000000000,
						cb8_1 = 32'b00001010001010000000000000000000,
						cb8_2 = 32'b00001010100011000000000000000000,
						cb8_3 = 32'b00001010111100000000000000000000,
						cb8_4 = 32'b00001011010101000000000000000000,
						cb8_5 = 32'b00001011101110000000000000000000,
						cb8_6 = 32'b00001100000111000000000000000000,
						cb8_7 = 32'b00001100100000000000000000000000,
						
						cb9_0 = 32'b00001011010101000000000000000000,
						cb9_1 = 32'b00001100000111000000000000000000,
						cb9_2 = 32'b00001100111001000000000000000000,
						cb9_3 = 32'b00001101101011000000000000000000;

//------------------------------------------------------------------
//                  -- State & Reg Declarations  --                   
//------------------------------------------------------------------

parameter START = 5'd0,
          INITVALUES = 5'd1,
          INITLOOP = 5'd2,
          CALCERROR = 5'd3,
			 POWERE = 5'd4,
          BESTECHECK = 5'd5,
          INCRJ = 5'd6,
          CHECKJ = 5'd7,
          CALCSE = 5'd8,
          DONE = 5'd9;

reg [3:0] STATE, NEXT_STATE;

//------------------------------------------------------------------
//                  -- Module Instantiations  --                   
//------------------------------------------------------------------

qadd #(Q,N) qadd0(cb0,{(vec[N-1] == 0)?1'b1:1'b0,vec[N-2:0]},out_e0); 		
qadd #(Q,N) qadd1(cb1,{(vec[N-1] == 0)?1'b1:1'b0,vec[N-2:0]},out_e1); 
qadd #(Q,N) qadd2(cb2,{(vec[N-1] == 0)?1'b1:1'b0,vec[N-2:0]},out_e2); 
qadd #(Q,N) qadd3(cb3,{(vec[N-1] == 0)?1'b1:1'b0,vec[N-2:0]},out_e3); 	
qadd #(Q,N) qadd4(cb4,{(vec[N-1] == 0)?1'b1:1'b0,vec[N-2:0]},out_e4); 
qadd #(Q,N) qadd5(cb5,{(vec[N-1] == 0)?1'b1:1'b0,vec[N-2:0]},out_e5); 
qadd #(Q,N) qadd6(cb6,{(vec[N-1] == 0)?1'b1:1'b0,vec[N-2:0]},out_e6); 
qadd #(Q,N) qadd7(cb7,{(vec[N-1] == 0)?1'b1:1'b0,vec[N-2:0]},out_e7); 
qadd #(Q,N) qadd8(cb8,{(vec[N-1] == 0)?1'b1:1'b0,vec[N-2:0]},out_e8); 
qadd #(Q,N) qadd9(cb9,{(vec[N-1] == 0)?1'b1:1'b0,vec[N-2:0]},out_e9); 
qadd #(Q,N) qadd10(cb10,{(vec[N-1] == 0)?1'b1:1'b0,vec[N-2:0]},out_e10); 
qadd #(Q,N) qadd11(cb11,{(vec[N-1] == 0)?1'b1:1'b0,vec[N-2:0]},out_e11); 
qadd #(Q,N) qadd12(cb12,{(vec[N-1] == 0)?1'b1:1'b0,vec[N-2:0]},out_e12); 
qadd #(Q,N) qadd13(cb13,{(vec[N-1] == 0)?1'b1:1'b0,vec[N-2:0]},out_e13); 
qadd #(Q,N) qadd14(cb14,{(vec[N-1] == 0)?1'b1:1'b0,vec[N-2:0]},out_e14); 
qadd #(Q,N) qadd15(cb15,{(vec[N-1] == 0)?1'b1:1'b0,vec[N-2:0]},out_e15); 	

fplessthan #(Q,N) fplt1(in_e,in_beste,lt1);

qmult #(Q,N) mult1(in_e1,in_e2,power_e);

//------------------------------------------------------------------
//                 -- Begin Declarations & Coding --                  
//------------------------------------------------------------------

always@(posedge clk or negedge rst)     // Determine STATE
begin

	if (rst == 1'b0)
		STATE <= START;
	else
		STATE <= NEXT_STATE;

end


always@(*)                              // Determine NEXT_STATE
begin
	case(STATE)

	START:
	begin
		if (startq) 
		begin
			NEXT_STATE = INITVALUES;
		end
		else
		begin
			NEXT_STATE = START;
		end
	end

	INITVALUES:
	begin
		NEXT_STATE = INITLOOP;
	end

	INITLOOP:
	begin
		NEXT_STATE = CALCERROR;
	end

	CALCERROR:
	begin
		NEXT_STATE = POWERE;
	end
	
	POWERE:
	begin
		NEXT_STATE = BESTECHECK;
	end

	BESTECHECK:
	begin
		NEXT_STATE = INCRJ;
	end

	INCRJ:
	begin
		NEXT_STATE = CHECKJ;
	end

	CHECKJ:
	begin
		if(j < m) 
		begin
			NEXT_STATE = INITLOOP;
		end
		else 
		begin
			NEXT_STATE = CALCSE;
		end
	end

	CALCSE:
	begin
		NEXT_STATE = DONE;
	end

	DONE:
	begin
		NEXT_STATE = START;
	end


	endcase
end


always@(posedge clk or negedge rst)     // Determine outputs
begin

	if (rst == 1'b0)
	begin
		besti <= 5'b0;
		e <= 32'b0;
		beste <= 32'b0_111111111111111_1111111111111111;
		j <= 5'd0;
		//startq <= 1'b0;
		doneq <= 1'b0;
	end

	else
	begin
		case(STATE)

		START:
		begin
			doneq <= 1'b0;
		end

		INITVALUES:
		begin
			besti <= 5'b0;
			beste <= 32'b0_111111111111111_1111111111111111;
			j <= 5'd0;
			//startq <= 1'b0;
		end

		INITLOOP:
		begin
			e <= 32'b0;
			case(orderi)
				5'd0: 
				begin
					cb0 <= cb0_0;
					cb1 <= cb0_1;
					cb2 <= cb0_2;
					cb3 <= cb0_3;
					cb4 <= cb0_4;
					cb5 <= cb0_5;
					cb6 <= cb0_6;
					cb7 <= cb0_7;
					cb8 <= cb0_8;
					cb9 <= cb0_9;
					cb10 <= cb0_10;
					cb11 <= cb0_11;
					cb12 <= cb0_12;
					cb13 <= cb0_13;
					cb14 <= cb0_14;
					cb15 <= cb0_15;
				end
				5'd1:
				begin
					cb0 <= cb1_0;
					cb1 <= cb1_1;
					cb2 <= cb1_2;
					cb3 <= cb1_3;
					cb4 <= cb1_4;
					cb5 <= cb1_5;
					cb6 <= cb1_6;
					cb7 <= cb1_7;
					cb8 <= cb1_8;
					cb9 <= cb1_9;
					cb10 <= cb1_10;
					cb11 <= cb1_11;
					cb12 <= cb1_12;
					cb13 <= cb1_13;
					cb14 <= cb1_14;
					cb15 <= cb1_15;
				end
				5'd2:
				begin
					cb0 <= cb2_0;
					cb1 <= cb2_1;
					cb2 <= cb2_2;
					cb3 <= cb2_3;
					cb4 <= cb2_4;
					cb5 <= cb2_5;
					cb6 <= cb2_6;
					cb7 <= cb2_7;
					cb8 <= cb2_8;
					cb9 <= cb2_9;
					cb10 <= cb2_10;
					cb11 <= cb2_11;
					cb12 <= cb2_12;
					cb13 <= cb2_13;
					cb14 <= cb2_14;
					cb15 <= cb2_15;
				end
				5'd3:
				begin
					cb0 <= cb3_0;
					cb1 <= cb3_1;
					cb2 <= cb3_2;
					cb3 <= cb3_3;
					cb4 <= cb3_4;
					cb5 <= cb3_5;
					cb6 <= cb3_6;
					cb7 <= cb3_7;
					cb8 <= cb3_8;
					cb9 <= cb3_9;
					cb10 <= cb3_10;
					cb11 <= cb3_11;
					cb12 <= cb3_12;
					cb13 <= cb3_13;
					cb14 <= cb3_14;
					cb15 <= cb3_15;
				end
				5'd4:
				begin
					cb0 <= cb4_0;
					cb1 <= cb4_1;
					cb2 <= cb4_2;
					cb3 <= cb4_3;
					cb4 <= cb4_4;
					cb5 <= cb4_5;
					cb6 <= cb4_6;
					cb7 <= cb4_7;
					cb8 <= cb4_8;
					cb9 <= cb4_9;
					cb10 <= cb4_10;
					cb11 <= cb4_11;
					cb12 <= cb4_12;
					cb13 <= cb4_13;
					cb14 <= cb4_14;
					cb15 <= cb4_15;
				end
				5'd5:
				begin
					cb0 <= cb5_0;
					cb1 <= cb5_1;
					cb2 <= cb5_2;
					cb3 <= cb5_3;
					cb4 <= cb5_4;
					cb5 <= cb5_5;
					cb6 <= cb5_6;
					cb7 <= cb5_7;
					cb8 <= cb5_8;
					cb9 <= cb5_9;
					cb10 <= cb5_10;
					cb11 <= cb5_11;
					cb12 <= cb5_12;
					cb13 <= cb5_13;
					cb14 <= cb5_14;
					cb15 <= cb5_15;
				end
				5'd6:
				begin
					cb0 <= cb6_0;
					cb1 <= cb6_1;
					cb2 <= cb6_2;
					cb3 <= cb6_3;
					cb4 <= cb6_4;
					cb5 <= cb6_5;
					cb6 <= cb6_6;
					cb7 <= cb6_7;
					cb8 <= cb6_8;
					cb9 <= cb6_9;
					cb10 <= cb6_10;
					cb11 <= cb6_11;
					cb12 <= cb6_12;
					cb13 <= cb6_13;
					cb14 <= cb6_14;
					cb15 <= cb6_15;
				end
				5'd7:
				begin
					cb0 <= cb7_0;
					cb1 <= cb7_1;
					cb2 <= cb7_2;
					cb3 <= cb7_3;
					cb4 <= cb7_4;
					cb5 <= cb7_5;
					cb6 <= cb7_6;
					cb7 <= cb7_7;
				end
				5'd8:
				begin
					cb0 <= cb8_0;
					cb1 <= cb8_1;
					cb2 <= cb8_2;
					cb3 <= cb8_3;
					cb4 <= cb8_4;
					cb5 <= cb8_5;
					cb6 <= cb8_6;
					cb7 <= cb8_7;
				end
				5'd9:
				begin
					cb0 <= cb9_0;
					cb1 <= cb9_1;
					cb2 <= cb9_2;
					cb3 <= cb9_3;
				end	
			endcase
		end

		CALCERROR:
		begin
			case(orderi)
				5'd0,5'd1,5'd2,5'd3,5'd4,5'd5,5'd6:
				begin
					case(j)
						5'd0: e <= out_e0;
						5'd1: e <= out_e1;
						5'd2: e <= out_e2;
						5'd3: e <= out_e3;
						5'd4: e <= out_e4;
						5'd5: e <= out_e5;
						5'd6: e <= out_e6;
						5'd7: e <= out_e7;
						5'd8: e <= out_e8;
						5'd9: e <= out_e9;
						5'd10: e <= out_e10;
						5'd11: e <= out_e11;
						5'd12: e <= out_e12;
						5'd13: e <= out_e13;
						5'd14: e <= out_e14;
						5'd15: e <= out_e15;
					endcase
				end
				5'd7,5'd8:
				begin
					case(j)
						5'd0: e <= out_e0;
						5'd1: e <= out_e1;
						5'd2: e <= out_e2;
						5'd3: e <= out_e3;
						5'd4: e <= out_e4;
						5'd5: e <= out_e5;
						5'd6: e <= out_e6;
						5'd7: e <= out_e7;
					endcase
				end
				5'd9:
				begin
					case(j)
						5'd0: e <= out_e0;
						5'd1: e <= out_e1;
						5'd2: e <= out_e2;
						5'd3: e <= out_e3;
					endcase
				end
			endcase
		end
		
		POWERE:
		begin
				in_e1 <= e;
				in_e2 <= e;
				abs_e <= {(e[N-1] == 1)?1'b0:1'b0,e[N-2:0]};
					 
				
		end

		BESTECHECK:
		begin
				in_e <= abs_e;
				in_beste <= beste;
				
			//	in_e <= 32'b1;
			//	in_beste <= 32'b111;
		end

		INCRJ:
		begin
				j <= j + 5'd1;
				if(lt1)
				begin
					beste <= abs_e;
					besti <= j;
				end
		end

		CHECKJ:
		begin
				
		end

		CALCSE:
		begin
			
		end

		DONE:
		begin
			doneq <= 1'b1;
		end

		endcase
	end

end


endmodule