/*
* Module         - ROM_cb6
* Top module     - cbselect
* Project        - CODEC2_ENCODE_2400
* Developer      - Santhiya S
* Date           - Mon Feb 04 15:19:31 2019
*
* Description    -
* Inputs         -
*static const float codes6[] = {
1500,
  1600,
  1700,
  1800,
  1900,
  2000,
  2100,
  2200,
  2300,
  2400,
  2500,
  2600,
  2700,
  2800,
  2900,
  3000
*};
*32 bits fixed point representation
   S - E  - M
   1 - 15 - 16
*/
module ROM_cb6(addr,dataout);

	parameter N = 32;
	input [3:0] addr;
	output reg [N-1:0] dataout;

	reg [N-1:0] cb6[15:0];
	
	always@(*)
	begin
			cb6[0] = 32'b00000101110111000000000000000000;
			cb6[1] = 32'b00000110010000000000000000000000;
			cb6[2] = 32'b00000110101001000000000000000000;
			cb6[3] = 32'b00000111000010000000000000000000;
			cb6[4] = 32'b00000111011011000000000000000000;
			cb6[5] = 32'b00000111110100000000000000000000;
			cb6[6] = 32'b00001000001101000000000000000000;
			cb6[7] = 32'b00001000100110000000000000000000;
			cb6[8] = 32'b00001000111111000000000000000000;
			cb6[9] = 32'b00001001011000000000000000000000;
			cb6[10] = 32'b00001001110001000000000000000000;
			cb6[11] = 32'b00001010001010000000000000000000;
			cb6[12] = 32'b00001010100011000000000000000000;
			cb6[13] = 32'b00001010111100000000000000000000;
			cb6[14] = 32'b00001011010101000000000000000000;
			cb6[15] = 32'b00001011101110000000000000000000;
		
		dataout = cb6[addr];
	end
endmodule
