/*
* Module         - ROM_nlp_fir[
* Top module     - cbselect
* Project        - CODEC2_ENCODE_2400
* Developer      - Santhiya S
* Date           - Mon Feb 04 15:19:31 2019
*
* Description    -
* Inputs         -

*32 bits fixed point representation
   S - E  - M
   1 - 15 - 16
*/
module ROM_nlp_fir(addr,dataout);

	parameter N = 80;
	input [5:0] addr;
	output reg [N-1:0] dataout;

	reg [N-1:0] nlp_fir[47:0];
	
	always@(*)
	begin
nlp_fir[0]  = 80'b10000000000000000000000000000000000000000000000000000000000000000000000001000110;
nlp_fir[1]  = 80'b10000000000000000000000000000000000000000000000000000000000000000000000001001000;
nlp_fir[2]  = 80'b10000000000000000000000000000000000000000000000000000000000000000000000000111100;
nlp_fir[3]  = 80'b10000000000000000000000000000000000000000000000000000000000000000000000000011011;
nlp_fir[4]  = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000100100;
nlp_fir[5]  = 80'b00000000000000000000000000000000000000000000000000000000000000000000000010000011;
nlp_fir[6]  = 80'b00000000000000000000000000000000000000000000000000000000000000000000000011110010;
nlp_fir[7]  = 80'b00000000000000000000000000000000000000000000000000000000000000000000000101010001;
nlp_fir[8]  = 80'b00000000000000000000000000000000000000000000000000000000000000000000000101101110;
nlp_fir[9]  = 80'b00000000000000000000000000000000000000000000000000000000000000000000000100011010;
nlp_fir[10]  = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000110100;
nlp_fir[11]  = 80'b10000000000000000000000000000000000000000000000000000000000000000000000100111011;
nlp_fir[12]  = 80'b10000000000000000000000000000000000000000000000000000000000000000000001011111111;
nlp_fir[13]  = 80'b10000000000000000000000000000000000000000000000000000000000000000000010010101000;
nlp_fir[14]  = 80'b10000000000000000000000000000000000000000000000000000000000000000000010110100110;
nlp_fir[15]  = 80'b10000000000000000000000000000000000000000000000000000000000000000000010101011011;
nlp_fir[16]  = 80'b10000000000000000000000000000000000000000000000000000000000000000000001101000111;
nlp_fir[17]  = 80'b00000000000000000000000000000000000000000000000000000000000000000000000011010011;
nlp_fir[18]  = 80'b00000000000000000000000000000000000000000000000000000000000000000000011011010100;
nlp_fir[19]  = 80'b00000000000000000000000000000000000000000000000000000000000000000000111000110110;
nlp_fir[20]  = 80'b00000000000000000000000000000000000000000000000000000000000000000001011000011000;
nlp_fir[21]  = 80'b00000000000000000000000000000000000000000000000000000000000000000001110101100011;
nlp_fir[22]  = 80'b00000000000000000000000000000000000000000000000000000000000000000010001100000001;
nlp_fir[23]  = 80'b00000000000000000000000000000000000000000000000000000000000000000010011000001111;
nlp_fir[24]  = 80'b00000000000000000000000000000000000000000000000000000000000000000010011000001111;
nlp_fir[25]  = 80'b00000000000000000000000000000000000000000000000000000000000000000010001100000001;
nlp_fir[26]  = 80'b00000000000000000000000000000000000000000000000000000000000000000001110101100011;
nlp_fir[27]  = 80'b00000000000000000000000000000000000000000000000000000000000000000001011000011000;
nlp_fir[28]  = 80'b00000000000000000000000000000000000000000000000000000000000000000000111000110110;
nlp_fir[29]  = 80'b00000000000000000000000000000000000000000000000000000000000000000000011011010100;
nlp_fir[30]  = 80'b00000000000000000000000000000000000000000000000000000000000000000000000011010011;
nlp_fir[31]  = 80'b10000000000000000000000000000000000000000000000000000000000000000000001101000111;
nlp_fir[32]  = 80'b10000000000000000000000000000000000000000000000000000000000000000000010101011011;
nlp_fir[33]  = 80'b10000000000000000000000000000000000000000000000000000000000000000000010110100110;
nlp_fir[34]  = 80'b10000000000000000000000000000000000000000000000000000000000000000000010010101000;
nlp_fir[35]  = 80'b10000000000000000000000000000000000000000000000000000000000000000000001011111111;
nlp_fir[36]  = 80'b10000000000000000000000000000000000000000000000000000000000000000000000100111011;
nlp_fir[37]  = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000110100;
nlp_fir[38]  = 80'b00000000000000000000000000000000000000000000000000000000000000000000000100011010;
nlp_fir[39]  = 80'b00000000000000000000000000000000000000000000000000000000000000000000000101101110;
nlp_fir[40]  = 80'b00000000000000000000000000000000000000000000000000000000000000000000000101010001;
nlp_fir[41]  = 80'b00000000000000000000000000000000000000000000000000000000000000000000000011110010;
nlp_fir[42]  = 80'b00000000000000000000000000000000000000000000000000000000000000000000000010000011;
nlp_fir[43]  = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000100100;
nlp_fir[44]  = 80'b10000000000000000000000000000000000000000000000000000000000000000000000000011011;
nlp_fir[45]  = 80'b10000000000000000000000000000000000000000000000000000000000000000000000000111100;
nlp_fir[46]  = 80'b10000000000000000000000000000000000000000000000000000000000000000000000001001000;
nlp_fir[47]  = 80'b10000000000000000000000000000000000000000000000000000000000000000000000001000110;
		
		dataout = nlp_fir[addr];
	end
endmodule
