/*
* Module         - find_nearest_weighted
* Top module     - encode_WoE
* Project        - CODEC2_ENCODE_2400
* Developer      - Santhiya S
* Date           - Thu Feb 07 14:48:10 2019
*
* Description    - 
* Inputs         - startfnw, x0,x1,w0,w1
* Simulation     - Waveform 24.vwf
*32 bits fixed point representation
   S - E  - M
   1 - 15 - 16
*/


module find_nearest_weighted (startfnw,clk,rst,x0,x1,w0,w1,nearest,donefnw);


//------------------------------------------------------------------
//                 -- Input/Output Declarations --                  
//------------------------------------------------------------------

	parameter N = 32;
	parameter Q = 16;
	
	input startfnw;
	input clk,rst;
	input [N-1:0] x0,x1,w0,w1;
	
	output reg [8:0] nearest;
	output reg donefnw;
	

//------------------------------------------------------------------
//                  -- State & Reg Declarations  --                   
//------------------------------------------------------------------

parameter START = 3'd0,
          INITVALUES = 3'd1,
          INITLOOP = 3'd2,
          CALCDIST = 3'd3,
          SETDIST = 3'd4,
          INCRI = 3'd5,
          CHECKI = 3'd6,
          DONE = 3'd7;

reg [2:0]STATE, NEXT_STATE;

//------------------------------------------------------------------
//                  -- Constants Declarations  --                   
//------------------------------------------------------------------

parameter [8:0] ndim = 9'd256; 

parameter [N-1:0] 	cb0 = 32'b00000000000000101011010111000010,
						cb1 = 32'b00000000000011000000010010110101,
						cb2 = 32'b00000000000000000000101111110111,
						cb3 = 32'b10000000000000101011110100100010,
						cb4 = 32'b00000000000000000001111011111001,
						cb5 = 32'b00000000000010000110001110010010,
						cb6 = 32'b10000000000000011001010010001101,
						cb7 = 32'b10000000000000001110010001101110,
						cb8 = 32'b00000000000000010011000101101101,
						cb9 = 32'b10000000000000011110101001100101,
						cb10 = 32'b00000000000000000010111111100101,
						cb11 = 32'b10000000000000110100011011011011,
						cb12 = 32'b00000000000000000101010100001110,
						cb13 = 32'b10000000000001111010101000011111,
						cb14 = 32'b10000000000000010111101010111100,
						cb15 = 32'b00000000000111110011111100000000,
						cb16 = 32'b00000000000000011000011100010001,
						cb17 = 32'b00000000000110111011010110100001,
						cb18 = 32'b10000000000000001000011000111101,
						cb19 = 32'b00000000000001010100000000000111,
						cb20 = 32'b00000000000000001000110110100111,
						cb21 = 32'b00000000000001110111000001010101,
						cb22 = 32'b10000000000000001101011111101100,
						cb23 = 32'b10000000000000011111001111110111,
						cb24 = 32'b00000000000000100100001110001110,
						cb25 = 32'b00000000000010001001110000111011,
						cb26 = 32'b00000000000000000010010010100101,
						cb27 = 32'b00000000000000100101110110010000,
						cb28 = 32'b00000000000000001001110111010011,
						cb29 = 32'b00000000000000010100100011000101,
						cb30 = 32'b10000000000000011011011000011001,
						cb31 = 32'b00000000000101100001100011000001,
						cb32 = 32'b00000000000000010000001000010100,
						cb33 = 32'b00000000000100010110010110000001,
						cb34 = 32'b10000000000000000001101101010001,
						cb35 = 32'b00000000000000010110101100111101,
						cb36 = 32'b10000000000000000010001011100001,
						cb37 = 32'b00000000000011100100011000001010,
						cb38 = 32'b10000000000000011011010110000110,
						cb39 = 32'b10000000000101001000100000101010,
						cb40 = 32'b00000000000000011010100001101010,
						cb41 = 32'b10000000000000110110010000011101,
						cb42 = 32'b00000000000000000010001101010111,
						cb43 = 32'b10000000000001001111010100110101,
						cb44 = 32'b00000000000000001000100101100111,
						cb45 = 32'b10000000000000011111000110011001,
						cb46 = 32'b00000000000000000011001001000001,
						cb47 = 32'b00000000001001001101101000010110,
						cb48 = 32'b00000000000000010100010111000001,
						cb49 = 32'b00000000000101101000111001110110,
						cb50 = 32'b10000000000000001010101110010011,
						cb51 = 32'b10000000000000011110011111110010,
						cb52 = 32'b00000000000000000110000111010000,
						cb53 = 32'b00000000000001100110011010110000,
						cb54 = 32'b10000000000000001100000111000100,
						cb55 = 32'b10000000000001001110011010101001,
						cb56 = 32'b00000000000000011101010001001101,
						cb57 = 32'b00000000000001001001110100100001,
						cb58 = 32'b00000000000000000101000110011100,
						cb59 = 32'b00000000000000001011110010100000,
						cb60 = 32'b00000000000000001001110011100001,
						cb61 = 32'b10000000000000100001001100110110,
						cb62 = 32'b10000000000000000110100011111111,
						cb63 = 32'b00000000000110001100100101111111,
						cb64 = 32'b00000000000000011100011010101001,
						cb65 = 32'b00000000000011010011000011011110,
						cb66 = 32'b00000000000000000001101101000000,
						cb67 = 32'b10000000000000000001101010111111,
						cb68 = 32'b00000000000000000011000100110100,
						cb69 = 32'b00000000000010100010111100001101,
						cb70 = 32'b10000000000000011101001100001101,
						cb71 = 32'b10000000000001111011011100110100,
						cb72 = 32'b00000000000000001110111001101100,
						cb73 = 32'b00000000000001000101100100101101,
						cb74 = 32'b00000000000000000100111100001110,
						cb75 = 32'b10000000000001000001011000000100,
						cb76 = 32'b00000000000000000110010110101011,
						cb77 = 32'b10000000000010111100111100010100,
						cb78 = 32'b10000000000000000000110001111000,
						cb79 = 32'b00000000001010010011101000110000,
						cb80 = 32'b00000000000000001110000010011001,
						cb81 = 32'b00000000001000111101100110101101,
						cb82 = 32'b10000000000000001100001010000001,
						cb83 = 32'b00000000000000000111101000000100,
						cb84 = 32'b00000000000000001111101010000101,
						cb85 = 32'b00000000000001111010110010110111,
						cb86 = 32'b10000000000000010011000111101111,
						cb87 = 32'b00000000000000110000100111110000,
						cb88 = 32'b00000000000000101010001111001111,
						cb89 = 32'b10000000000000110110100100111011,
						cb90 = 32'b00000000000000000011000011101101,
						cb91 = 32'b00000000000000111001101001111111,
						cb92 = 32'b00000000000000000110011100100110,
						cb93 = 32'b00000000000000010001010110010100,
						cb94 = 32'b10000000000000100010011011101010,
						cb95 = 32'b00000000000100100001101110001011,
						cb96 = 32'b00000000000000011000101111111011,
						cb97 = 32'b00000000000010000101001010011101,
						cb98 = 32'b10000000000000000010010010100001,
						cb99 = 32'b10000000000001000001001101101111,
						cb100 = 32'b10000000000000000010011001101111,
						cb101 = 32'b00000000000001011101110111100010,
						cb102 = 32'b10000000000000010110100010001111,
						cb103 = 32'b10000000000000110100000000101101,
						cb104 = 32'b00000000000000011001000011101111,
						cb105 = 32'b10000000000010100110100111000111,
						cb106 = 32'b00000000000000000010110110011100,
						cb107 = 32'b10000000000010100011101000001001,
						cb108 = 32'b00000000000000000101110010110110,
						cb109 = 32'b10000000000000000000011101001111,
						cb110 = 32'b10000000000000000001000111110011,
						cb111 = 32'b00000000000110000110010000000100,
						cb112 = 32'b00000000000000001001100001000001,
						cb113 = 32'b00000000000100010111101110011000,
						cb114 = 32'b10000000000000000100100101110111,
						cb115 = 32'b10000000000001101110011101110001,
						cb116 = 32'b00000000000000000111011011111110,
						cb117 = 32'b00000000000010100011010010011011,
						cb118 = 32'b10000000000000010000000111000000,
						cb119 = 32'b10000000000011100101101101110001,
						cb120 = 32'b00000000000000100101010001011110,
						cb121 = 32'b10000000000000111011000100001101,
						cb122 = 32'b00000000000000000101010111110011,
						cb123 = 32'b00000000000000100110100000111010,
						cb124 = 32'b00000000000000010000010100001000,
						cb125 = 32'b10000000000000110010011111011000,
						cb126 = 32'b10000000000000010100001001101011,
						cb127 = 32'b00000000000001111111110111101101,
						cb128 = 32'b00000000000000100110001000111001,
						cb129 = 32'b00000000000100111010111000111011,
						cb130 = 32'b10000000000000000001100001001110,
						cb131 = 32'b10000000000000100110100111101010,
						cb132 = 32'b00000000000000000011010110010110,
						cb133 = 32'b00000000000001101010101000101110,
						cb134 = 32'b10000000000000100011100010010101,
						cb135 = 32'b00000000000000010110000100111110,
						cb136 = 32'b00000000000000010100101011011010,
						cb137 = 32'b00000000000000100000101111011100,
						cb138 = 32'b00000000000000000011111001011110,
						cb139 = 32'b10000000000000001110010000000111,
						cb140 = 32'b00000000000000000110110111000100,
						cb141 = 32'b10000000000001110011000110010011,
						cb142 = 32'b10000000000000010001110100011110,
						cb143 = 32'b00000000001010010101011101100101,
						cb144 = 32'b00000000000000101001110000011011,
						cb145 = 32'b00000000000111110010001111110111,
						cb146 = 32'b10000000000000000111001001001011,
						cb147 = 32'b00000000000000101000100011000000,
						cb148 = 32'b00000000000000000111110101110111,
						cb149 = 32'b00000000000001001010000010101000,
						cb150 = 32'b10000000000000010001111000000010,
						cb151 = 32'b10000000000000110011110111100010,
						cb152 = 32'b00000000000000011100101010100011,
						cb153 = 32'b00000000000010000110101000111000,
						cb154 = 32'b00000000000000000010011111110000,
						cb155 = 32'b00000000000000000010111011101111,
						cb156 = 32'b00000000000000001000100001001110,
						cb157 = 32'b00000000000000110010011110010000,
						cb158 = 32'b10000000000000001100001110110101,
						cb159 = 32'b00000000000100101000001110010101,
						cb160 = 32'b00000000000000001111001111010000,
						cb161 = 32'b00000000000010111100010101110011,
						cb162 = 32'b10000000000000000101010100100011,
						cb163 = 32'b00000000000000000101100011010100,
						cb164 = 32'b00000000000000000011001111000001,
						cb165 = 32'b00000000000011101011011110000000,
						cb166 = 32'b10000000000000100010000100010101,
						cb167 = 32'b10000000000011111000111100011010,
						cb168 = 32'b00000000000000010101101010000100,
						cb169 = 32'b10000000000000011110110101000010,
						cb170 = 32'b10000000000000000000001011001110,
						cb171 = 32'b10000000000100000101011000011110,
						cb172 = 32'b00000000000000000110011000101000,
						cb173 = 32'b10000000000000101100101001100010,
						cb174 = 32'b00000000000000001100000000101011,
						cb175 = 32'b00000000000111110010010111110110,
						cb176 = 32'b00000000000000001010011111011110,
						cb177 = 32'b00000000000110000111101101011101,
						cb178 = 32'b10000000000000000111010000000101,
						cb179 = 32'b10000000000000001011110001100010,
						cb180 = 32'b00000000000000000100100101110010,
						cb181 = 32'b00000000000001101000101111110100,
						cb182 = 32'b10000000000000001011011100110110,
						cb183 = 32'b10000000000011000101101110011000,
						cb184 = 32'b00000000000000011000110001101001,
						cb185 = 32'b00000000000000111101111101000110,
						cb186 = 32'b00000000000000000100010110011001,
						cb187 = 32'b00000000000000001100110101100110,
						cb188 = 32'b00000000000000001000000010000111,
						cb189 = 32'b10000000000001001101101011010111,
						cb190 = 32'b10000000000000000111111100111101,
						cb191 = 32'b00000000000100011100001100001011,
						cb192 = 32'b00000000000000010011000011101111,
						cb193 = 32'b00000000000011011111010001010011,
						cb194 = 32'b00000000000000000000010000000000,
						cb195 = 32'b00000000000000010101010011100001,
						cb196 = 32'b00000000000000000101011110000100,
						cb197 = 32'b00000000000010001110111101110100,
						cb198 = 32'b10000000000000100101000011100110,
						cb199 = 32'b10000000000001010110010100100010,
						cb200 = 32'b00000000000000001100001000110100,
						cb201 = 32'b00000000000000011111011011101001,
						cb202 = 32'b00000000000000000011110111000111,
						cb203 = 32'b10000000000000110011110011011001,
						cb204 = 32'b00000000000000000100010001100100,
						cb205 = 32'b10000000000010110011110000000001,
						cb206 = 32'b10000000000000000100010111101011,
						cb207 = 32'b00000000001000001001111111110010,
						cb208 = 32'b00000000000000011100000011100110,
						cb209 = 32'b00000000001010000110111010010111,
						cb210 = 32'b10000000000000001100100010110100,
						cb211 = 32'b00000000000000110000101110110110,
						cb212 = 32'b00000000000000001011010010111011,
						cb213 = 32'b00000000000001011010100101000011,
						cb214 = 32'b10000000000000010110001011101011,
						cb215 = 32'b00000000000000010101101010000010,
						cb216 = 32'b00000000000000100110000001011111,
						cb217 = 32'b00000000000000011010110011000010,
						cb218 = 32'b00000000000000000011111000110011,
						cb219 = 32'b00000000000001001011101101110000,
						cb220 = 32'b00000000000000000111110111000001,
						cb221 = 32'b00000000000000000101101010100011,
						cb222 = 32'b10000000000000011001101101010100,
						cb223 = 32'b00000000000010001010100010110000,
						cb224 = 32'b00000000000000010010101011000111,
						cb225 = 32'b00000000000001011111110010110010,
						cb226 = 32'b10000000000000000010001100111001,
						cb227 = 32'b10000000000011000000101010101100,
						cb228 = 32'b10000000000000000100000001011010,
						cb229 = 32'b00000000000010100110010110101110,
						cb230 = 32'b10000000000000010110111001110111,
						cb231 = 32'b10000000000010001110011101110011,
						cb232 = 32'b00000000000000001111110011111111,
						cb233 = 32'b10000000000011010011010110000001,
						cb234 = 32'b00000000000000000100001011110000,
						cb235 = 32'b10000000000001100101101011011111,
						cb236 = 32'b00000000000000000110010101011011,
						cb237 = 32'b10000000000000001011001111011000,
						cb238 = 32'b00000000000000000100100010100000,
						cb239 = 32'b00000000000110101110011001001100,
						cb240 = 32'b00000000000000000110101111000011,
						cb241 = 32'b00000000000011110111000100011001,
						cb242 = 32'b10000000000000000101101100010101,
						cb243 = 32'b10000000000011011011101001010001,
						cb244 = 32'b00000000000000001000011100000001,
						cb245 = 32'b00000000000011000110011000000100,
						cb246 = 32'b10000000000000010010101101101000,
						cb247 = 32'b10000000000011111111111110011101,
						cb248 = 32'b00000000000000011110100000011100,
						cb249 = 32'b10000000000001011101000011101000,
						cb250 = 32'b00000000000000000101101010111111,
						cb251 = 32'b00000000000000111101101000000000,
						cb252 = 32'b00000000000000001101001101100101,
						cb253 = 32'b10000000000001000010100110100010,
						cb254 = 32'b10000000000000000111110101111101,
						cb255 = 32'b00000000000011010000111010100100,
						cb256 = 32'b00000000000000100100000101111010,
						cb257 = 32'b00000000000011011000011011000010,
						cb258 = 32'b10000000000000000000000101000100,
						cb259 = 32'b10000000000000110011110010110100,
						cb260 = 32'b00000000000000000000011011010110,
						cb261 = 32'b00000000000001111101110111001111,
						cb262 = 32'b10000000000000011100111101110100,
						cb263 = 32'b10000000000000000111001110000000,
						cb264 = 32'b00000000000000010001010101110101,
						cb265 = 32'b10000000000000000010111100000001,
						cb266 = 32'b00000000000000000010001011000110,
						cb267 = 32'b10000000000000100100010000111110,
						cb268 = 32'b00000000000000000110000000110101,
						cb269 = 32'b10000000000001011000001100100010,
						cb270 = 32'b10000000000000011111011101101000,
						cb271 = 32'b00000000001001101010111011010010,
						cb272 = 32'b00000000000000011111101001011101,
						cb273 = 32'b00000000000110001001000011000100,
						cb274 = 32'b10000000000000001011010001100100,
						cb275 = 32'b00000000000001100101101111011010,
						cb276 = 32'b00000000000000000111101100010100,
						cb277 = 32'b00000000000001110000110100111111,
						cb278 = 32'b10000000000000001111100111110110,
						cb279 = 32'b10000000000000100110110000111000,
						cb280 = 32'b00000000000000101000000010001100,
						cb281 = 32'b00000000000001101100001001100100,
						cb282 = 32'b00000000000000000001010101100110,
						cb283 = 32'b00000000000000110100001001000000,
						cb284 = 32'b00000000000000001000101100101011,
						cb285 = 32'b00000000000000001110100011110110,
						cb286 = 32'b10000000000000010011101101100001,
						cb287 = 32'b00000000000101110001011101101100,
						cb288 = 32'b00000000000000001100100100010110,
						cb289 = 32'b00000000000011101100111010010111,
						cb290 = 32'b10000000000000000011011010101011,
						cb291 = 32'b00000000000000011011000000100000,
						cb292 = 32'b00000000000000000000000100110111,
						cb293 = 32'b00000000000100100010101111111011,
						cb294 = 32'b10000000000000011000110000010100,
						cb295 = 32'b10000000000100000001110111100110,
						cb296 = 32'b00000000000000011000000001000100,
						cb297 = 32'b10000000000000110100011111111000,
						cb298 = 32'b00000000000000000001010010000011,
						cb299 = 32'b10000000000001001010001001111101,
						cb300 = 32'b00000000000000000111101000000001,
						cb301 = 32'b10000000000000100010111001010001,
						cb302 = 32'b00000000000000000111000101000101,
						cb303 = 32'b00000000001010000100110111010010,
						cb304 = 32'b00000000000000010001001010100001,
						cb305 = 32'b00000000000110111001011110001101,
						cb306 = 32'b10000000000000001001100001000000,
						cb307 = 32'b10000000000001000010101010110100,
						cb308 = 32'b00000000000000000110110000100111,
						cb309 = 32'b00000000000001111001110110111000,
						cb310 = 32'b10000000000000001110110101110010,
						cb311 = 32'b10000000000001110100011000111111,
						cb312 = 32'b00000000000000011111110111011010,
						cb313 = 32'b00000000000000010100101111011110,
						cb314 = 32'b00000000000000000100101010010011,
						cb315 = 32'b00000000000000100110011000010110,
						cb316 = 32'b00000000000000001011100010011000,
						cb317 = 32'b10000000000000011111001101011011,
						cb318 = 32'b10000000000000001100110111100011,
						cb319 = 32'b00000000000110001110110111110011,
						cb320 = 32'b00000000000000011010010111111100,
						cb321 = 32'b00000000000100110001111010100100,
						cb322 = 32'b00000000000000000000111110010011,
						cb323 = 32'b10000000000000001001011100110100,
						cb324 = 32'b00000000000000000100010000011110,
						cb325 = 32'b00000000000010010001101001101110,
						cb326 = 32'b10000000000000011111010100011000,
						cb327 = 32'b10000000000000101110001001110101,
						cb328 = 32'b00000000000000010001110111101111,
						cb329 = 32'b00000000000000101010110000100010,
						cb330 = 32'b00000000000000000101101011000101,
						cb331 = 32'b10000000000000101011111110100000,
						cb332 = 32'b00000000000000000101010010101010,
						cb333 = 32'b10000000000011100010011111110110,
						cb334 = 32'b10000000000000001000011100100001,
						cb335 = 32'b00000000001001111001001101011010,
						cb336 = 32'b00000000000000001111110110111100,
						cb337 = 32'b00000000001010110011000111101011,
						cb338 = 32'b10000000000000001001011011110001,
						cb339 = 32'b00000000000000010100010011101001,
						cb340 = 32'b00000000000000001100100110010011,
						cb341 = 32'b00000000000010001011101100001111,
						cb342 = 32'b10000000000000010000001110001000,
						cb343 = 32'b00000000000000010000011001101010,
						cb344 = 32'b00000000000000101101001101001101,
						cb345 = 32'b00000000000000011110010100110111,
						cb346 = 32'b00000000000000000011110110101010,
						cb347 = 32'b00000000000000101011111011011101,
						cb348 = 32'b00000000000000000110110101011100,
						cb349 = 32'b00000000000000101000101101100001,
						cb350 = 32'b10000000000000011111001111111111,
						cb351 = 32'b00000000000011000011111001110110,
						cb352 = 32'b00000000000000010111001011011000,
						cb353 = 32'b00000000000011000000111110001010,
						cb354 = 32'b10000000000000000011010111100010,
						cb355 = 32'b10000000000000110110000100001010,
						cb356 = 32'b10000000000000000000111010000100,
						cb357 = 32'b00000000000010100011010000111001,
						cb358 = 32'b10000000000000011010011100000001,
						cb359 = 32'b10000000000001010001101001001101,
						cb360 = 32'b00000000000000010100101101110100,
						cb361 = 32'b10000000000011000100010101010011,
						cb362 = 32'b00000000000000000001110010010010,
						cb363 = 32'b10000000000010001010110100001001,
						cb364 = 32'b00000000000000000101001110011110,
						cb365 = 32'b10000000000000010010101011101001,
						cb366 = 32'b00000000000000000000010110010011,
						cb367 = 32'b00000000000111110010000000110100,
						cb368 = 32'b00000000000000000111010010010000,
						cb369 = 32'b00000000000101010111011111101001,
						cb370 = 32'b10000000000000000110000000011100,
						cb371 = 32'b10000000000000110101111100000111,
						cb372 = 32'b00000000000000000110010011000100,
						cb373 = 32'b00000000000010110100110101001111,
						cb374 = 32'b10000000000000001101100111111001,
						cb375 = 32'b10000000000100110110101000110110,
						cb376 = 32'b00000000000000100001101101100110,
						cb377 = 32'b10000000000000100011101010010110,
						cb378 = 32'b00000000000000000101111110001100,
						cb379 = 32'b00000000000000011110110010001111,
						cb380 = 32'b00000000000000001110001001101010,
						cb381 = 32'b10000000000000011011100001110111,
						cb382 = 32'b10000000000000001111100110100001,
						cb383 = 32'b00000000000010011101011100010010,
						cb384 = 32'b00000000000000100000000011011000,
						cb385 = 32'b00000000000100010110010100111000,
						cb386 = 32'b10000000000000000000100101110011,
						cb387 = 32'b10000000000000010001110010000010,
						cb388 = 32'b00000000000000000010011000000001,
						cb389 = 32'b00000000000001010110011001100100,
						cb390 = 32'b10000000000000011110101000010110,
						cb391 = 32'b00000000000001001100011000011001,
						cb392 = 32'b00000000000000010111001010101010,
						cb393 = 32'b00000000000000001000100110000000,
						cb394 = 32'b00000000000000000011000111101010,
						cb395 = 32'b10000000000000010000100111000110,
						cb396 = 32'b00000000000000000111111011101010,
						cb397 = 32'b10000000000010011111010001111100,
						cb398 = 32'b10000000000000010000111100011001,
						cb399 = 32'b00000000001000001111001001110101,
						cb400 = 32'b00000000000000100000001011011111,
						cb401 = 32'b00000000001000000111010001010011,
						cb402 = 32'b10000000000000000100111101000101,
						cb403 = 32'b00000000000001001011100000010111,
						cb404 = 32'b00000000000000000110111110100011,
						cb405 = 32'b00000000000001001010001010110001,
						cb406 = 32'b10000000000000010011110010110011,
						cb407 = 32'b10000000000000010100000100011000,
						cb408 = 32'b00000000000000100000010111010010,
						cb409 = 32'b00000000000010010110110110100111,
						cb410 = 32'b00000000000000000011000010111010,
						cb411 = 32'b00000000000000010111010111110101,
						cb412 = 32'b00000000000000000111101010100000,
						cb413 = 32'b00000000000000100111110000011011,
						cb414 = 32'b10000000000000010001010000010111,
						cb415 = 32'b00000000000100000011100011000001,
						cb416 = 32'b00000000000000010011010100100111,
						cb417 = 32'b00000000000010011010011101111010,
						cb418 = 32'b10000000000000000100001000010001,
						cb419 = 32'b10000000000000011010110000011111,
						cb420 = 32'b00000000000000000001001001100100,
						cb421 = 32'b00000000000011010110101001111110,
						cb422 = 32'b10000000000000011110000010010010,
						cb423 = 32'b10000000000100000001001001101110,
						cb424 = 32'b00000000000000010100101000100001,
						cb425 = 32'b10000000000001001101111100000101,
						cb426 = 32'b00000000000000000001000101010101,
						cb427 = 32'b10000000000011010111000101010100,
						cb428 = 32'b00000000000000000110111110000000,
						cb429 = 32'b10000000000001000010101001011110,
						cb430 = 32'b00000000000000000111011101010100,
						cb431 = 32'b00000000000111101001011011101001,
						cb432 = 32'b00000000000000001110011110100111,
						cb433 = 32'b00000000000101011001100100010110,
						cb434 = 32'b10000000000000001000010010110011,
						cb435 = 32'b10000000000000101000100000110100,
						cb436 = 32'b00000000000000000101011001011101,
						cb437 = 32'b00000000000001011010001100100011,
						cb438 = 32'b10000000000000001000111000010010,
						cb439 = 32'b10000000000100010110011010000111,
						cb440 = 32'b00000000000000011011000100011111,
						cb441 = 32'b00000000000000010010010101001111,
						cb442 = 32'b00000000000000000011101001011001,
						cb443 = 32'b00000000000000001110001110101000,
						cb444 = 32'b00000000000000001001011001011001,
						cb445 = 32'b10000000000001011011101011001111,
						cb446 = 32'b10000000000000000100001100011011,
						cb447 = 32'b00000000000100101010101010100110,
						cb448 = 32'b00000000000000010110010100100001,
						cb449 = 32'b00000000000100010000000010111110,
						cb450 = 32'b10000000000000000000010011100011,
						cb451 = 32'b00000000000001000100111011110001,
						cb452 = 32'b00000000000000000100110111100010,
						cb453 = 32'b00000000000011001010101101111110,
						cb454 = 32'b10000000000000100001001011110101,
						cb455 = 32'b10000000000001100111010111111001,
						cb456 = 32'b00000000000000001110101110101000,
						cb457 = 32'b00000000000000010011011010000100,
						cb458 = 32'b00000000000000000100100011110000,
						cb459 = 32'b10000000000000011100100100010100,
						cb460 = 32'b00000000000000000011010110110000,
						cb461 = 32'b10000000000100000000011000100100,
						cb462 = 32'b10000000000000001010001011010101,
						cb463 = 32'b00000000000111111001001110101001,
						cb464 = 32'b00000000000000010101100110010010,
						cb465 = 32'b00000000001000101010110101110000,
						cb466 = 32'b10000000000000001111100010111100,
						cb467 = 32'b00000000000001010100110100000101,
						cb468 = 32'b00000000000000001001011100011010,
						cb469 = 32'b00000000000001000111001100100000,
						cb470 = 32'b10000000000000011001000101011111,
						cb471 = 32'b00000000000000111001101000110110,
						cb472 = 32'b00000000000000100010010100111111,
						cb473 = 32'b00000000000001001000010001000011,
						cb474 = 32'b00000000000000000100101111001000,
						cb475 = 32'b00000000000001000001111011000011,
						cb476 = 32'b00000000000000000111000111111111,
						cb477 = 32'b00000000000000001101111001100111,
						cb478 = 32'b10000000000000010111000100100010,
						cb479 = 32'b00000000000011100010000011011110,
						cb480 = 32'b00000000000000010101101100010010,
						cb481 = 32'b00000000000001100000000111100100,
						cb482 = 32'b10000000000000000000001101000111,
						cb483 = 32'b10000000000001110111111100011111,
						cb484 = 32'b10000000000000000110111000010100,
						cb485 = 32'b00000000000010001000000000000111,
						cb486 = 32'b10000000000000010011010001100110,
						cb487 = 32'b10000000000001110001110011111110,
						cb488 = 32'b00000000000000010001100111011100,
						cb489 = 32'b10000000000001101101011000111001,
						cb490 = 32'b00000000000000000011001001001011,
						cb491 = 32'b10000000000001100011101111100111,
						cb492 = 32'b00000000000000000110111111001110,
						cb493 = 32'b10000000000000010010000100111001,
						cb494 = 32'b00000000000000000010010000011011,
						cb495 = 32'b00000000000101101101101011011010,
						cb496 = 32'b00000000000000000100101001110011,
						cb497 = 32'b00000000000100101100111110110111,
						cb498 = 32'b10000000000000001000011110001111,
						cb499 = 32'b10000000000001111011101110000101,
						cb500 = 32'b00000000000000001010001001100000,
						cb501 = 32'b00000000000010101100101000110000,
						cb502 = 32'b10000000000000010101010110110000,
						cb503 = 32'b10000000000101000101001101100111,
						cb504 = 32'b00000000000000011101000011001101,
						cb505 = 32'b10000000000000011110011100111111,
						cb506 = 32'b00000000000000000110010100010000,
						cb507 = 32'b00000000000000111100110000101110,
						cb508 = 32'b00000000000000001011101110010001,
						cb509 = 32'b10000000000010000010111100001110,
						cb510 = 32'b10000000000000001011110111000010,
						cb511 = 32'b00000000000010111100010010101111;


//------------------------------------------------------------------
//                  -- Module Instatntiations  --                   
//------------------------------------------------------------------

wire lt1;
reg [8:0] i;
reg [N-1:0] in_cb0,in_cb1,distance,min_dist,comp1,comp2;
wire [N-1:0] xcb0,xcb1,sq_xcb0,sq_xcb1,out_dist0,out_dist1,
				 out_dist;
				 
reg [N-1:0]  dist0, dist1;
				 

qadd #(Q,N) adder1(x0,{(in_cb0[N-1] == 0)?1'b1:1'b0,in_cb0[N-2:0]},xcb0);
qadd #(Q,N) adder2(x1,{(in_cb1[N-1] == 0)?1'b1:1'b0,in_cb1[N-2:0]},xcb1);

qmult #(Q,N) mult1(xcb0,xcb0,sq_xcb0);
qmult #(Q,N) mult2(xcb1,xcb1,sq_xcb1);
qmult #(Q,N) mult3(w0,sq_xcb0,out_dist0);
qmult #(Q,N) mult4(w1,sq_xcb1,out_dist1);

qadd #(Q,N) adder3(dist0,dist1,out_dist);

fplessthan #(Q,N) fplt1(comp1,comp2,lt1);



//------------------------------------------------------------------
//                 -- Begin Declarations & Coding --                  
//------------------------------------------------------------------

always@(posedge clk or negedge rst)     // Determine STATE
begin

	if (rst == 1'b0)
		STATE <= START;
	else
		STATE <= NEXT_STATE;

end


always@(*)                              // Determine NEXT_STATE
begin
	case(STATE)

	START:
	begin
		if(startfnw == 1'b1)
		begin
			NEXT_STATE = INITVALUES;
		end
		else
		begin
			NEXT_STATE = START;
		end
	end

	INITVALUES:
	begin
		NEXT_STATE = INITLOOP;
	end

	INITLOOP:
	begin
		NEXT_STATE = CALCDIST;
	end

	CALCDIST:
	begin
		NEXT_STATE = SETDIST;
	end

	SETDIST:
	begin
		NEXT_STATE = INCRI;
	end

	INCRI:
	begin
		NEXT_STATE = CHECKI;
	end

	CHECKI:
	begin
		if(i < ndim)
		begin
			NEXT_STATE = INITLOOP;
		end
		else
		begin
			NEXT_STATE = DONE;
		end
	end

	DONE:
	begin
		NEXT_STATE = START;
	end

	endcase
end


always@(posedge clk or negedge rst)     // Determine outputs
begin

	if (rst == 1'b0)
	begin
		donefnw <= 1'b0;
		nearest <= 9'b0;
		i <= 9'b0;
	end

	else
	begin
		case(STATE)

		START:
		begin
			donefnw <= 1'b0;
		end

		INITVALUES:
		begin
			min_dist <= 32'b01111111111111111111111111111111;
			nearest <= 9'b0;
			i <= 9'b0;
		end

		INITLOOP:
		begin
			distance <= 32'b0;
			case (i)
			9'd0:
			begin
				in_cb0 <= cb0;
				in_cb1 <= cb1;
			end
			9'd1:
			begin
				in_cb0 <= cb2;
				in_cb1 <= cb3;
			end
			9'd2:
			begin
				in_cb0 <= cb4;
				in_cb1 <= cb5;
			end
			9'd3:
			begin
				in_cb0 <= cb6;
				in_cb1 <= cb7;
			end
			9'd4:
			begin
				in_cb0 <= cb8;
				in_cb1 <= cb9;
			end
			9'd5:
			begin
				in_cb0 <= cb10;
				in_cb1 <= cb11;
			end
			9'd6:
			begin
				in_cb0 <= cb12;
				in_cb1 <= cb13;
			end
			9'd7:
			begin
				in_cb0 <= cb14;
				in_cb1 <= cb15;
			end
			9'd8:
			begin
				in_cb0 <= cb16;
				in_cb1 <= cb17;
			end
			9'd9:
			begin
				in_cb0 <= cb18;
				in_cb1 <= cb19;
			end
			9'd10:
			begin
				in_cb0 <= cb20;
				in_cb1 <= cb21;
			end
			9'd11:
			begin
				in_cb0 <= cb22;
				in_cb1 <= cb23;
			end
			9'd12:
			begin
				in_cb0 <= cb24;
				in_cb1 <= cb25;
			end
			9'd13:
			begin
				in_cb0 <= cb26;
				in_cb1 <= cb27;
			end
			9'd14:
			begin
				in_cb0 <= cb28;
				in_cb1 <= cb29;
			end
			9'd15:
			begin
				in_cb0 <= cb30;
				in_cb1 <= cb31;
			end
			9'd16:
			begin
				in_cb0 <= cb32;
				in_cb1 <= cb33;
			end
			9'd17:
			begin
				in_cb0 <= cb34;
				in_cb1 <= cb35;
			end
			9'd18:
			begin
				in_cb0 <= cb36;
				in_cb1 <= cb37;
			end
			9'd19:
			begin
				in_cb0 <= cb38;
				in_cb1 <= cb39;
			end
			9'd20:
			begin
				in_cb0 <= cb40;
				in_cb1 <= cb41;
			end
			9'd21:
			begin
				in_cb0 <= cb42;
				in_cb1 <= cb43;
			end
			9'd22:
			begin
				in_cb0 <= cb44;
				in_cb1 <= cb45;
			end
			9'd23:
			begin
				in_cb0 <= cb46;
				in_cb1 <= cb47;
			end
			9'd24:
			begin
				in_cb0 <= cb48;
				in_cb1 <= cb49;
			end
			9'd25:
			begin
				in_cb0 <= cb50;
				in_cb1 <= cb51;
			end
			9'd26:
			begin
				in_cb0 <= cb52;
				in_cb1 <= cb53;
			end
			9'd27:
			begin
				in_cb0 <= cb54;
				in_cb1 <= cb55;
			end
			9'd28:
			begin
				in_cb0 <= cb56;
				in_cb1 <= cb57;
			end
			9'd29:
			begin
				in_cb0 <= cb58;
				in_cb1 <= cb59;
			end
			9'd30:
			begin
				in_cb0 <= cb60;
				in_cb1 <= cb61;
			end
			9'd31:
			begin
				in_cb0 <= cb62;
				in_cb1 <= cb63;
			end
			9'd32:
			begin
				in_cb0 <= cb64;
				in_cb1 <= cb65;
			end
			9'd33:
			begin
				in_cb0 <= cb66;
				in_cb1 <= cb67;
			end
			9'd34:
			begin
				in_cb0 <= cb68;
				in_cb1 <= cb69;
			end
			9'd35:
			begin
				in_cb0 <= cb70;
				in_cb1 <= cb71;
			end
			9'd36:
			begin
				in_cb0 <= cb72;
				in_cb1 <= cb73;
			end
			9'd37:
			begin
				in_cb0 <= cb74;
				in_cb1 <= cb75;
			end
			9'd38:
			begin
				in_cb0 <= cb76;
				in_cb1 <= cb77;
			end
			9'd39:
			begin
				in_cb0 <= cb78;
				in_cb1 <= cb79;
			end
			9'd40:
			begin
				in_cb0 <= cb80;
				in_cb1 <= cb81;
			end
			9'd41:
			begin
				in_cb0 <= cb82;
				in_cb1 <= cb83;
			end
			9'd42:
			begin
				in_cb0 <= cb84;
				in_cb1 <= cb85;
			end
			9'd43:
			begin
				in_cb0 <= cb86;
				in_cb1 <= cb87;
			end
			9'd44:
			begin
				in_cb0 <= cb88;
				in_cb1 <= cb89;
			end
			9'd45:
			begin
				in_cb0 <= cb90;
				in_cb1 <= cb91;
			end
			9'd46:
			begin
				in_cb0 <= cb92;
				in_cb1 <= cb93;
			end
			9'd47:
			begin
				in_cb0 <= cb94;
				in_cb1 <= cb95;
			end
			9'd48:
			begin
				in_cb0 <= cb96;
				in_cb1 <= cb97;
			end
			9'd49:
			begin
				in_cb0 <= cb98;
				in_cb1 <= cb99;
			end
			9'd50:
			begin
				in_cb0 <= cb100;
				in_cb1 <= cb101;
			end
			9'd51:
			begin
				in_cb0 <= cb102;
				in_cb1 <= cb103;
			end
			9'd52:
			begin
				in_cb0 <= cb104;
				in_cb1 <= cb105;
			end
			9'd53:
			begin
				in_cb0 <= cb106;
				in_cb1 <= cb107;
			end
			9'd54:
			begin
				in_cb0 <= cb108;
				in_cb1 <= cb109;
			end
			9'd55:
			begin
				in_cb0 <= cb110;
				in_cb1 <= cb111;
			end
			9'd56:
			begin
				in_cb0 <= cb112;
				in_cb1 <= cb113;
			end
			9'd57:
			begin
				in_cb0 <= cb114;
				in_cb1 <= cb115;
			end
			9'd58:
			begin
				in_cb0 <= cb116;
				in_cb1 <= cb117;
			end
			9'd59:
			begin
				in_cb0 <= cb118;
				in_cb1 <= cb119;
			end
			9'd60:
			begin
				in_cb0 <= cb120;
				in_cb1 <= cb121;
			end
			9'd61:
			begin
				in_cb0 <= cb122;
				in_cb1 <= cb123;
			end
			9'd62:
			begin
				in_cb0 <= cb124;
				in_cb1 <= cb125;
			end
			9'd63:
			begin
				in_cb0 <= cb126;
				in_cb1 <= cb127;
			end
			9'd64:
			begin
				in_cb0 <= cb128;
				in_cb1 <= cb129;
			end
			9'd65:
			begin
				in_cb0 <= cb130;
				in_cb1 <= cb131;
			end
			9'd66:
			begin
				in_cb0 <= cb132;
				in_cb1 <= cb133;
			end
			9'd67:
			begin
				in_cb0 <= cb134;
				in_cb1 <= cb135;
			end
			9'd68:
			begin
				in_cb0 <= cb136;
				in_cb1 <= cb137;
			end
			9'd69:
			begin
				in_cb0 <= cb138;
				in_cb1 <= cb139;
			end
			9'd70:
			begin
				in_cb0 <= cb140;
				in_cb1 <= cb141;
			end
			9'd71:
			begin
				in_cb0 <= cb142;
				in_cb1 <= cb143;
			end
			9'd72:
			begin
				in_cb0 <= cb144;
				in_cb1 <= cb145;
			end
			9'd73:
			begin
				in_cb0 <= cb146;
				in_cb1 <= cb147;
			end
			9'd74:
			begin
				in_cb0 <= cb148;
				in_cb1 <= cb149;
			end
			9'd75:
			begin
				in_cb0 <= cb150;
				in_cb1 <= cb151;
			end
			9'd76:
			begin
				in_cb0 <= cb152;
				in_cb1 <= cb153;
			end
			9'd77:
			begin
				in_cb0 <= cb154;
				in_cb1 <= cb155;
			end
			9'd78:
			begin
				in_cb0 <= cb156;
				in_cb1 <= cb157;
			end
			9'd79:
			begin
				in_cb0 <= cb158;
				in_cb1 <= cb159;
			end
			9'd80:
			begin
				in_cb0 <= cb160;
				in_cb1 <= cb161;
			end
			9'd81:
			begin
				in_cb0 <= cb162;
				in_cb1 <= cb163;
			end
			9'd82:
			begin
				in_cb0 <= cb164;
				in_cb1 <= cb165;
			end
			9'd83:
			begin
				in_cb0 <= cb166;
				in_cb1 <= cb167;
			end
			9'd84:
			begin
				in_cb0 <= cb168;
				in_cb1 <= cb169;
			end
			9'd85:
			begin
				in_cb0 <= cb170;
				in_cb1 <= cb171;
			end
			9'd86:
			begin
				in_cb0 <= cb172;
				in_cb1 <= cb173;
			end
			9'd87:
			begin
				in_cb0 <= cb174;
				in_cb1 <= cb175;
			end
			9'd88:
			begin
				in_cb0 <= cb176;
				in_cb1 <= cb177;
			end
			9'd89:
			begin
				in_cb0 <= cb178;
				in_cb1 <= cb179;
			end
			9'd90:
			begin
				in_cb0 <= cb180;
				in_cb1 <= cb181;
			end
			9'd91:
			begin
				in_cb0 <= cb182;
				in_cb1 <= cb183;
			end
			9'd92:
			begin
				in_cb0 <= cb184;
				in_cb1 <= cb185;
			end
			9'd93:
			begin
				in_cb0 <= cb186;
				in_cb1 <= cb187;
			end
			9'd94:
			begin
				in_cb0 <= cb188;
				in_cb1 <= cb189;
			end
			9'd95:
			begin
				in_cb0 <= cb190;
				in_cb1 <= cb191;
			end
			9'd96:
			begin
				in_cb0 <= cb192;
				in_cb1 <= cb193;
			end
			9'd97:
			begin
				in_cb0 <= cb194;
				in_cb1 <= cb195;
			end
			9'd98:
			begin
				in_cb0 <= cb196;
				in_cb1 <= cb197;
			end
			9'd99:
			begin
				in_cb0 <= cb198;
				in_cb1 <= cb199;
			end
			9'd100:
			begin
				in_cb0 <= cb200;
				in_cb1 <= cb201;
			end
			9'd101:
			begin
				in_cb0 <= cb202;
				in_cb1 <= cb203;
			end
			9'd102:
			begin
				in_cb0 <= cb204;
				in_cb1 <= cb205;
			end
			9'd103:
			begin
				in_cb0 <= cb206;
				in_cb1 <= cb207;
			end
			9'd104:
			begin
				in_cb0 <= cb208;
				in_cb1 <= cb209;
			end
			9'd105:
			begin
				in_cb0 <= cb210;
				in_cb1 <= cb211;
			end
			9'd106:
			begin
				in_cb0 <= cb212;
				in_cb1 <= cb213;
			end
			9'd107:
			begin
				in_cb0 <= cb214;
				in_cb1 <= cb215;
			end
			9'd108:
			begin
				in_cb0 <= cb216;
				in_cb1 <= cb217;
			end
			9'd109:
			begin
				in_cb0 <= cb218;
				in_cb1 <= cb219;
			end
			9'd110:
			begin
				in_cb0 <= cb220;
				in_cb1 <= cb221;
			end
			9'd111:
			begin
				in_cb0 <= cb222;
				in_cb1 <= cb223;
			end
			9'd112:
			begin
				in_cb0 <= cb224;
				in_cb1 <= cb225;
			end
			9'd113:
			begin
				in_cb0 <= cb226;
				in_cb1 <= cb227;
			end
			9'd114:
			begin
				in_cb0 <= cb228;
				in_cb1 <= cb229;
			end
			9'd115:
			begin
				in_cb0 <= cb230;
				in_cb1 <= cb231;
			end
			9'd116:
			begin
				in_cb0 <= cb232;
				in_cb1 <= cb233;
			end
			9'd117:
			begin
				in_cb0 <= cb234;
				in_cb1 <= cb235;
			end
			9'd118:
			begin
				in_cb0 <= cb236;
				in_cb1 <= cb237;
			end
			9'd119:
			begin
				in_cb0 <= cb238;
				in_cb1 <= cb239;
			end
			9'd120:
			begin
				in_cb0 <= cb240;
				in_cb1 <= cb241;
			end
			9'd121:
			begin
				in_cb0 <= cb242;
				in_cb1 <= cb243;
			end
			9'd122:
			begin
				in_cb0 <= cb244;
				in_cb1 <= cb245;
			end
			9'd123:
			begin
				in_cb0 <= cb246;
				in_cb1 <= cb247;
			end
			9'd124:
			begin
				in_cb0 <= cb248;
				in_cb1 <= cb249;
			end
			9'd125:
			begin
				in_cb0 <= cb250;
				in_cb1 <= cb251;
			end
			9'd126:
			begin
				in_cb0 <= cb252;
				in_cb1 <= cb253;
			end
			9'd127:
			begin
				in_cb0 <= cb254;
				in_cb1 <= cb255;
			end
			9'd128:
			begin
				in_cb0 <= cb256;
				in_cb1 <= cb257;
			end
			9'd129:
			begin
				in_cb0 <= cb258;
				in_cb1 <= cb259;
			end
			9'd130:
			begin
				in_cb0 <= cb260;
				in_cb1 <= cb261;
			end
			9'd131:
			begin
				in_cb0 <= cb262;
				in_cb1 <= cb263;
			end
			9'd132:
			begin
				in_cb0 <= cb264;
				in_cb1 <= cb265;
			end
			9'd133:
			begin
				in_cb0 <= cb266;
				in_cb1 <= cb267;
			end
			9'd134:
			begin
				in_cb0 <= cb268;
				in_cb1 <= cb269;
			end
			9'd135:
			begin
				in_cb0 <= cb270;
				in_cb1 <= cb271;
			end
			9'd136:
			begin
				in_cb0 <= cb272;
				in_cb1 <= cb273;
			end
			9'd137:
			begin
				in_cb0 <= cb274;
				in_cb1 <= cb275;
			end
			9'd138:
			begin
				in_cb0 <= cb276;
				in_cb1 <= cb277;
			end
			9'd139:
			begin
				in_cb0 <= cb278;
				in_cb1 <= cb279;
			end
			9'd140:
			begin
				in_cb0 <= cb280;
				in_cb1 <= cb281;
			end
			9'd141:
			begin
				in_cb0 <= cb282;
				in_cb1 <= cb283;
			end
			9'd142:
			begin
				in_cb0 <= cb284;
				in_cb1 <= cb285;
			end
			9'd143:
			begin
				in_cb0 <= cb286;
				in_cb1 <= cb287;
			end
			9'd144:
			begin
				in_cb0 <= cb288;
				in_cb1 <= cb289;
			end
			9'd145:
			begin
				in_cb0 <= cb290;
				in_cb1 <= cb291;
			end
			9'd146:
			begin
				in_cb0 <= cb292;
				in_cb1 <= cb293;
			end
			9'd147:
			begin
				in_cb0 <= cb294;
				in_cb1 <= cb295;
			end
			9'd148:
			begin
				in_cb0 <= cb296;
				in_cb1 <= cb297;
			end
			9'd149:
			begin
				in_cb0 <= cb298;
				in_cb1 <= cb299;
			end
			9'd150:
			begin
				in_cb0 <= cb300;
				in_cb1 <= cb301;
			end
			9'd151:
			begin
				in_cb0 <= cb302;
				in_cb1 <= cb303;
			end
			9'd152:
			begin
				in_cb0 <= cb304;
				in_cb1 <= cb305;
			end
			9'd153:
			begin
				in_cb0 <= cb306;
				in_cb1 <= cb307;
			end
			9'd154:
			begin
				in_cb0 <= cb308;
				in_cb1 <= cb309;
			end
			9'd155:
			begin
				in_cb0 <= cb310;
				in_cb1 <= cb311;
			end
			9'd156:
			begin
				in_cb0 <= cb312;
				in_cb1 <= cb313;
			end
			9'd157:
			begin
				in_cb0 <= cb314;
				in_cb1 <= cb315;
			end
			9'd158:
			begin
				in_cb0 <= cb316;
				in_cb1 <= cb317;
			end
			9'd159:
			begin
				in_cb0 <= cb318;
				in_cb1 <= cb319;
			end
			9'd160:
			begin
				in_cb0 <= cb320;
				in_cb1 <= cb321;
			end
			9'd161:
			begin
				in_cb0 <= cb322;
				in_cb1 <= cb323;
			end
			9'd162:
			begin
				in_cb0 <= cb324;
				in_cb1 <= cb325;
			end
			9'd163:
			begin
				in_cb0 <= cb326;
				in_cb1 <= cb327;
			end
			9'd164:
			begin
				in_cb0 <= cb328;
				in_cb1 <= cb329;
			end
			9'd165:
			begin
				in_cb0 <= cb330;
				in_cb1 <= cb331;
			end
			9'd166:
			begin
				in_cb0 <= cb332;
				in_cb1 <= cb333;
			end
			9'd167:
			begin
				in_cb0 <= cb334;
				in_cb1 <= cb335;
			end
			9'd168:
			begin
				in_cb0 <= cb336;
				in_cb1 <= cb337;
			end
			9'd169:
			begin
				in_cb0 <= cb338;
				in_cb1 <= cb339;
			end
			9'd170:
			begin
				in_cb0 <= cb340;
				in_cb1 <= cb341;
			end
			9'd171:
			begin
				in_cb0 <= cb342;
				in_cb1 <= cb343;
			end
			9'd172:
			begin
				in_cb0 <= cb344;
				in_cb1 <= cb345;
			end
			9'd173:
			begin
				in_cb0 <= cb346;
				in_cb1 <= cb347;
			end
			9'd174:
			begin
				in_cb0 <= cb348;
				in_cb1 <= cb349;
			end
			9'd175:
			begin
				in_cb0 <= cb350;
				in_cb1 <= cb351;
			end
			9'd176:
			begin
				in_cb0 <= cb352;
				in_cb1 <= cb353;
			end
			9'd177:
			begin
				in_cb0 <= cb354;
				in_cb1 <= cb355;
			end
			9'd178:
			begin
				in_cb0 <= cb356;
				in_cb1 <= cb357;
			end
			9'd179:
			begin
				in_cb0 <= cb358;
				in_cb1 <= cb359;
			end
			9'd180:
			begin
				in_cb0 <= cb360;
				in_cb1 <= cb361;
			end
			9'd181:
			begin
				in_cb0 <= cb362;
				in_cb1 <= cb363;
			end
			9'd182:
			begin
				in_cb0 <= cb364;
				in_cb1 <= cb365;
			end
			9'd183:
			begin
				in_cb0 <= cb366;
				in_cb1 <= cb367;
			end
			9'd184:
			begin
				in_cb0 <= cb368;
				in_cb1 <= cb369;
			end
			9'd185:
			begin
				in_cb0 <= cb370;
				in_cb1 <= cb371;
			end
			9'd186:
			begin
				in_cb0 <= cb372;
				in_cb1 <= cb373;
			end
			9'd187:
			begin
				in_cb0 <= cb374;
				in_cb1 <= cb375;
			end
			9'd188:
			begin
				in_cb0 <= cb376;
				in_cb1 <= cb377;
			end
			9'd189:
			begin
				in_cb0 <= cb378;
				in_cb1 <= cb379;
			end
			9'd190:
			begin
				in_cb0 <= cb380;
				in_cb1 <= cb381;
			end
			9'd191:
			begin
				in_cb0 <= cb382;
				in_cb1 <= cb383;
			end
			9'd192:
			begin
				in_cb0 <= cb384;
				in_cb1 <= cb385;
			end
			9'd193:
			begin
				in_cb0 <= cb386;
				in_cb1 <= cb387;
			end
			9'd194:
			begin
				in_cb0 <= cb388;
				in_cb1 <= cb389;
			end
			9'd195:
			begin
				in_cb0 <= cb390;
				in_cb1 <= cb391;
			end
			9'd196:
			begin
				in_cb0 <= cb392;
				in_cb1 <= cb393;
			end
			9'd197:
			begin
				in_cb0 <= cb394;
				in_cb1 <= cb395;
			end
			9'd198:
			begin
				in_cb0 <= cb396;
				in_cb1 <= cb397;
			end
			9'd199:
			begin
				in_cb0 <= cb398;
				in_cb1 <= cb399;
			end
			9'd200:
			begin
				in_cb0 <= cb400;
				in_cb1 <= cb401;
			end
			9'd201:
			begin
				in_cb0 <= cb402;
				in_cb1 <= cb403;
			end
			9'd202:
			begin
				in_cb0 <= cb404;
				in_cb1 <= cb405;
			end
			9'd203:
			begin
				in_cb0 <= cb406;
				in_cb1 <= cb407;
			end
			9'd204:
			begin
				in_cb0 <= cb408;
				in_cb1 <= cb409;
			end
			9'd205:
			begin
				in_cb0 <= cb410;
				in_cb1 <= cb411;
			end
			9'd206:
			begin
				in_cb0 <= cb412;
				in_cb1 <= cb413;
			end
			9'd207:
			begin
				in_cb0 <= cb414;
				in_cb1 <= cb415;
			end
			9'd208:
			begin
				in_cb0 <= cb416;
				in_cb1 <= cb417;
			end
			9'd209:
			begin
				in_cb0 <= cb418;
				in_cb1 <= cb419;
			end
			9'd210:
			begin
				in_cb0 <= cb420;
				in_cb1 <= cb421;
			end
			9'd211:
			begin
				in_cb0 <= cb422;
				in_cb1 <= cb423;
			end
			9'd212:
			begin
				in_cb0 <= cb424;
				in_cb1 <= cb425;
			end
			9'd213:
			begin
				in_cb0 <= cb426;
				in_cb1 <= cb427;
			end
			9'd214:
			begin
				in_cb0 <= cb428;
				in_cb1 <= cb429;
			end
			9'd215:
			begin
				in_cb0 <= cb430;
				in_cb1 <= cb431;
			end
			9'd216:
			begin
				in_cb0 <= cb432;
				in_cb1 <= cb433;
			end
			9'd217:
			begin
				in_cb0 <= cb434;
				in_cb1 <= cb435;
			end
			9'd218:
			begin
				in_cb0 <= cb436;
				in_cb1 <= cb437;
			end
			9'd219:
			begin
				in_cb0 <= cb438;
				in_cb1 <= cb439;
			end
			9'd220:
			begin
				in_cb0 <= cb440;
				in_cb1 <= cb441;
			end
			9'd221:
			begin
				in_cb0 <= cb442;
				in_cb1 <= cb443;
			end
			9'd222:
			begin
				in_cb0 <= cb444;
				in_cb1 <= cb445;
			end
			9'd223:
			begin
				in_cb0 <= cb446;
				in_cb1 <= cb447;
			end
			9'd224:
			begin
				in_cb0 <= cb448;
				in_cb1 <= cb449;
			end
			9'd225:
			begin
				in_cb0 <= cb450;
				in_cb1 <= cb451;
			end
			9'd226:
			begin
				in_cb0 <= cb452;
				in_cb1 <= cb453;
			end
			9'd227:
			begin
				in_cb0 <= cb454;
				in_cb1 <= cb455;
			end
			9'd228:
			begin
				in_cb0 <= cb456;
				in_cb1 <= cb457;
			end
			9'd229:
			begin
				in_cb0 <= cb458;
				in_cb1 <= cb459;
			end
			9'd230:
			begin
				in_cb0 <= cb460;
				in_cb1 <= cb461;
			end
			9'd231:
			begin
				in_cb0 <= cb462;
				in_cb1 <= cb463;
			end
			9'd232:
			begin
				in_cb0 <= cb464;
				in_cb1 <= cb465;
			end
			9'd233:
			begin
				in_cb0 <= cb466;
				in_cb1 <= cb467;
			end
			9'd234:
			begin
				in_cb0 <= cb468;
				in_cb1 <= cb469;
			end
			9'd235:
			begin
				in_cb0 <= cb470;
				in_cb1 <= cb471;
			end
			9'd236:
			begin
				in_cb0 <= cb472;
				in_cb1 <= cb473;
			end
			9'd237:
			begin
				in_cb0 <= cb474;
				in_cb1 <= cb475;
			end
			9'd238:
			begin
				in_cb0 <= cb476;
				in_cb1 <= cb477;
			end
			9'd239:
			begin
				in_cb0 <= cb478;
				in_cb1 <= cb479;
			end
			9'd240:
			begin
				in_cb0 <= cb480;
				in_cb1 <= cb481;
			end
			9'd241:
			begin
				in_cb0 <= cb482;
				in_cb1 <= cb483;
			end
			9'd242:
			begin
				in_cb0 <= cb484;
				in_cb1 <= cb485;
			end
			9'd243:
			begin
				in_cb0 <= cb486;
				in_cb1 <= cb487;
			end
			9'd244:
			begin
				in_cb0 <= cb488;
				in_cb1 <= cb489;
			end
			9'd245:
			begin
				in_cb0 <= cb490;
				in_cb1 <= cb491;
			end
			9'd246:
			begin
				in_cb0 <= cb492;
				in_cb1 <= cb493;
			end
			9'd247:
			begin
				in_cb0 <= cb494;
				in_cb1 <= cb495;
			end
			9'd248:
			begin
				in_cb0 <= cb496;
				in_cb1 <= cb497;
			end
			9'd249:
			begin
				in_cb0 <= cb498;
				in_cb1 <= cb499;
			end
			9'd250:
			begin
				in_cb0 <= cb500;
				in_cb1 <= cb501;
			end
			9'd251:
			begin
				in_cb0 <= cb502;
				in_cb1 <= cb503;
			end
			9'd252:
			begin
				in_cb0 <= cb504;
				in_cb1 <= cb505;
			end
			9'd253:
			begin
				in_cb0 <= cb506;
				in_cb1 <= cb507;
			end
			9'd254:
			begin
				in_cb0 <= cb508;
				in_cb1 <= cb509;
			end
			9'd255:
			begin
				in_cb0 <= cb510;
				in_cb1 <= cb511;
			end
			endcase
			
		end

		CALCDIST:
		begin
			dist0 <= out_dist0;
			dist1 <= out_dist1;
		end

		SETDIST:
		begin
			distance <= out_dist;
			comp1 <= out_dist;
			comp2 <= min_dist;
		end

		INCRI:
		begin
			i <= i + 9'd1;
			if(lt1)
			begin
				min_dist <= distance;
				nearest <= i;
			end
		end

		CHECKI:
		begin
			
		end

		DONE:
		begin
			donefnw <= 1'b1;
		end

		endcase
	end
	end

endmodule