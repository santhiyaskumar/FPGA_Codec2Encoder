/*
* Module         - ROM_speech_w[[
* Top module     - cbselect
* Project        - CODEC2_ENCODE_2400
* Developer      - Santhiya S
* Date           - Mon Feb 04 15:19:31 2019
*
* Description    -
* Inputs         -

*32 bits fixed point representation
   S - E  - M
   1 - 15 - 16
*/
module ROM_speech_w(addr,dataout);

	parameter N = 32;
	input [9:0] addr;
	output reg [N-1:0] dataout;

	reg [N-1:0] w[319:0];
	
	always@(*)
	begin

					w[0]  = 32'b00000000000000000000000000000000;
					w[1]  = 32'b00000000000000000000000000000000;
					w[2]  = 32'b00000000000000000000000000000000;
					w[3]  = 32'b00000000000000000000000000000000;
					w[4]  = 32'b00000000000000000000000000000000;
					w[5]  = 32'b00000000000000000000000000000000;
					w[6]  = 32'b00000000000000000000000000000000;
					w[7]  = 32'b00000000000000000000000000000000;
					w[8]  = 32'b00000000000000000000000000000000;
					w[9]  = 32'b00000000000000000000000000000000;
					w[10]  = 32'b00000000000000000000000000000000;
					w[11]  = 32'b00000000000000000000000000000000;
					w[12]  = 32'b00000000000000000000000000000000;
					w[13]  = 32'b00000000000000000000000000000000;
					w[14]  = 32'b00000000000000000000000000000000;
					w[15]  = 32'b00000000000000000000000000000000;
					w[16]  = 32'b00000000000000000000000000000000;
					w[17]  = 32'b00000000000000000000000000000000;
					w[18]  = 32'b00000000000000000000000000000000;
					w[19]  = 32'b00000000000000000000000000000000;
					w[20]  = 32'b00000000000000000000000000000000;
					w[21]  = 32'b00000000000000000000000000000000;
					w[22]  = 32'b00000000000000000000000000000000;
					w[23]  = 32'b00000000000000000000000000000000;
					w[24]  = 32'b00000000000000000000000000000000;
					w[25]  = 32'b00000000000000000000000000000000;
					w[26]  = 32'b00000000000000000000000000000000;
					w[27]  = 32'b00000000000000000000000000000001;
					w[28]  = 32'b00000000000000000000000000000001;
					w[29]  = 32'b00000000000000000000000000000010;
					w[30]  = 32'b00000000000000000000000000000010;
					w[31]  = 32'b00000000000000000000000000000011;
					w[32]  = 32'b00000000000000000000000000000100;
					w[33]  = 32'b00000000000000000000000000000101;
					w[34]  = 32'b00000000000000000000000000000110;
					w[35]  = 32'b00000000000000000000000000000111;
					w[36]  = 32'b00000000000000000000000000001000;
					w[37]  = 32'b00000000000000000000000000001001;
					w[38]  = 32'b00000000000000000000000000001010;
					w[39]  = 32'b00000000000000000000000000001011;
					w[40]  = 32'b00000000000000000000000000001100;
					w[41]  = 32'b00000000000000000000000000001110;
					w[42]  = 32'b00000000000000000000000000001111;
					w[43]  = 32'b00000000000000000000000000010001;
					w[44]  = 32'b00000000000000000000000000010010;
					w[45]  = 32'b00000000000000000000000000010100;
					w[46]  = 32'b00000000000000000000000000010110;
					w[47]  = 32'b00000000000000000000000000010111;
					w[48]  = 32'b00000000000000000000000000011001;
					w[49]  = 32'b00000000000000000000000000011011;
					w[50]  = 32'b00000000000000000000000000011101;
					w[51]  = 32'b00000000000000000000000000011111;
					w[52]  = 32'b00000000000000000000000000100001;
					w[53]  = 32'b00000000000000000000000000100011;
					w[54]  = 32'b00000000000000000000000000100101;
					w[55]  = 32'b00000000000000000000000000100111;
					w[56]  = 32'b00000000000000000000000000101010;
					w[57]  = 32'b00000000000000000000000000101100;
					w[58]  = 32'b00000000000000000000000000101110;
					w[59]  = 32'b00000000000000000000000000110001;
					w[60]  = 32'b00000000000000000000000000110011;
					w[61]  = 32'b00000000000000000000000000110110;
					w[62]  = 32'b00000000000000000000000000111000;
					w[63]  = 32'b00000000000000000000000000111011;
					w[64]  = 32'b00000000000000000000000000111101;
					w[65]  = 32'b00000000000000000000000001000000;
					w[66]  = 32'b00000000000000000000000001000011;
					w[67]  = 32'b00000000000000000000000001000101;
					w[68]  = 32'b00000000000000000000000001001000;
					w[69]  = 32'b00000000000000000000000001001011;
					w[70]  = 32'b00000000000000000000000001001110;
					w[71]  = 32'b00000000000000000000000001010001;
					w[72]  = 32'b00000000000000000000000001010100;
					w[73]  = 32'b00000000000000000000000001010111;
					w[74]  = 32'b00000000000000000000000001011010;
					w[75]  = 32'b00000000000000000000000001011101;
					w[76]  = 32'b00000000000000000000000001100000;
					w[77]  = 32'b00000000000000000000000001100011;
					w[78]  = 32'b00000000000000000000000001100110;
					w[79]  = 32'b00000000000000000000000001101001;
					w[80]  = 32'b00000000000000000000000001101100;
					w[81]  = 32'b00000000000000000000000001101111;
					w[82]  = 32'b00000000000000000000000001110010;
					w[83]  = 32'b00000000000000000000000001110101;
					w[84]  = 32'b00000000000000000000000001111001;
					w[85]  = 32'b00000000000000000000000001111100;
					w[86]  = 32'b00000000000000000000000001111111;
					w[87]  = 32'b00000000000000000000000010000010;
					w[88]  = 32'b00000000000000000000000010000101;
					w[89]  = 32'b00000000000000000000000010001001;
					w[90]  = 32'b00000000000000000000000010001100;
					w[91]  = 32'b00000000000000000000000010001111;
					w[92]  = 32'b00000000000000000000000010010010;
					w[93]  = 32'b00000000000000000000000010010101;
					w[94]  = 32'b00000000000000000000000010011001;
					w[95]  = 32'b00000000000000000000000010011100;
					w[96]  = 32'b00000000000000000000000010011111;
					w[97]  = 32'b00000000000000000000000010100010;
					w[98]  = 32'b00000000000000000000000010100101;
					w[99]  = 32'b00000000000000000000000010101000;
					w[100]  = 32'b00000000000000000000000010101100;
					w[101]  = 32'b00000000000000000000000010101111;
					w[102]  = 32'b00000000000000000000000010110010;
					w[103]  = 32'b00000000000000000000000010110101;
					w[104]  = 32'b00000000000000000000000010111000;
					w[105]  = 32'b00000000000000000000000010111011;
					w[106]  = 32'b00000000000000000000000010111110;
					w[107]  = 32'b00000000000000000000000011000001;
					w[108]  = 32'b00000000000000000000000011000100;
					w[109]  = 32'b00000000000000000000000011000111;
					w[110]  = 32'b00000000000000000000000011001010;
					w[111]  = 32'b00000000000000000000000011001101;
					w[112]  = 32'b00000000000000000000000011010000;
					w[113]  = 32'b00000000000000000000000011010010;
					w[114]  = 32'b00000000000000000000000011010101;
					w[115]  = 32'b00000000000000000000000011011000;
					w[116]  = 32'b00000000000000000000000011011011;
					w[117]  = 32'b00000000000000000000000011011101;
					w[118]  = 32'b00000000000000000000000011100000;
					w[119]  = 32'b00000000000000000000000011100011;
					w[120]  = 32'b00000000000000000000000011100101;
					w[121]  = 32'b00000000000000000000000011101000;
					w[122]  = 32'b00000000000000000000000011101010;
					w[123]  = 32'b00000000000000000000000011101100;
					w[124]  = 32'b00000000000000000000000011101111;
					w[125]  = 32'b00000000000000000000000011110001;
					w[126]  = 32'b00000000000000000000000011110011;
					w[127]  = 32'b00000000000000000000000011110110;
					w[128]  = 32'b00000000000000000000000011111000;
					w[129]  = 32'b00000000000000000000000011111010;
					w[130]  = 32'b00000000000000000000000011111100;
					w[131]  = 32'b00000000000000000000000011111110;
					w[132]  = 32'b00000000000000000000000100000000;
					w[133]  = 32'b00000000000000000000000100000010;
					w[134]  = 32'b00000000000000000000000100000011;
					w[135]  = 32'b00000000000000000000000100000101;
					w[136]  = 32'b00000000000000000000000100000111;
					w[137]  = 32'b00000000000000000000000100001000;
					w[138]  = 32'b00000000000000000000000100001010;
					w[139]  = 32'b00000000000000000000000100001011;
					w[140]  = 32'b00000000000000000000000100001101;
					w[141]  = 32'b00000000000000000000000100001110;
					w[142]  = 32'b00000000000000000000000100010000;
					w[143]  = 32'b00000000000000000000000100010001;
					w[144]  = 32'b00000000000000000000000100010010;
					w[145]  = 32'b00000000000000000000000100010011;
					w[146]  = 32'b00000000000000000000000100010100;
					w[147]  = 32'b00000000000000000000000100010101;
					w[148]  = 32'b00000000000000000000000100010110;
					w[149]  = 32'b00000000000000000000000100010111;
					w[150]  = 32'b00000000000000000000000100011000;
					w[151]  = 32'b00000000000000000000000100011000;
					w[152]  = 32'b00000000000000000000000100011001;
					w[153]  = 32'b00000000000000000000000100011001;
					w[154]  = 32'b00000000000000000000000100011010;
					w[155]  = 32'b00000000000000000000000100011010;
					w[156]  = 32'b00000000000000000000000100011011;
					w[157]  = 32'b00000000000000000000000100011011;
					w[158]  = 32'b00000000000000000000000100011011;
					w[159]  = 32'b00000000000000000000000100011011;
					w[160]  = 32'b00000000000000000000000100011011;
					w[161]  = 32'b00000000000000000000000100011011;
					w[162]  = 32'b00000000000000000000000100011011;
					w[163]  = 32'b00000000000000000000000100011011;
					w[164]  = 32'b00000000000000000000000100011011;
					w[165]  = 32'b00000000000000000000000100011010;
					w[166]  = 32'b00000000000000000000000100011010;
					w[167]  = 32'b00000000000000000000000100011001;
					w[168]  = 32'b00000000000000000000000100011001;
					w[169]  = 32'b00000000000000000000000100011000;
					w[170]  = 32'b00000000000000000000000100011000;
					w[171]  = 32'b00000000000000000000000100010111;
					w[172]  = 32'b00000000000000000000000100010110;
					w[173]  = 32'b00000000000000000000000100010101;
					w[174]  = 32'b00000000000000000000000100010100;
					w[175]  = 32'b00000000000000000000000100010011;
					w[176]  = 32'b00000000000000000000000100010010;
					w[177]  = 32'b00000000000000000000000100010001;
					w[178]  = 32'b00000000000000000000000100010000;
					w[179]  = 32'b00000000000000000000000100001110;
					w[180]  = 32'b00000000000000000000000100001101;
					w[181]  = 32'b00000000000000000000000100001011;
					w[182]  = 32'b00000000000000000000000100001010;
					w[183]  = 32'b00000000000000000000000100001000;
					w[184]  = 32'b00000000000000000000000100000111;
					w[185]  = 32'b00000000000000000000000100000101;
					w[186]  = 32'b00000000000000000000000100000011;
					w[187]  = 32'b00000000000000000000000100000010;
					w[188]  = 32'b00000000000000000000000100000000;
					w[189]  = 32'b00000000000000000000000011111110;
					w[190]  = 32'b00000000000000000000000011111100;
					w[191]  = 32'b00000000000000000000000011111010;
					w[192]  = 32'b00000000000000000000000011111000;
					w[193]  = 32'b00000000000000000000000011110110;
					w[194]  = 32'b00000000000000000000000011110011;
					w[195]  = 32'b00000000000000000000000011110001;
					w[196]  = 32'b00000000000000000000000011101111;
					w[197]  = 32'b00000000000000000000000011101100;
					w[198]  = 32'b00000000000000000000000011101010;
					w[199]  = 32'b00000000000000000000000011101000;
					w[200]  = 32'b00000000000000000000000011100101;
					w[201]  = 32'b00000000000000000000000011100011;
					w[202]  = 32'b00000000000000000000000011100000;
					w[203]  = 32'b00000000000000000000000011011101;
					w[204]  = 32'b00000000000000000000000011011011;
					w[205]  = 32'b00000000000000000000000011011000;
					w[206]  = 32'b00000000000000000000000011010101;
					w[207]  = 32'b00000000000000000000000011010010;
					w[208]  = 32'b00000000000000000000000011010000;
					w[209]  = 32'b00000000000000000000000011001101;
					w[210]  = 32'b00000000000000000000000011001010;
					w[211]  = 32'b00000000000000000000000011000111;
					w[212]  = 32'b00000000000000000000000011000100;
					w[213]  = 32'b00000000000000000000000011000001;
					w[214]  = 32'b00000000000000000000000010111110;
					w[215]  = 32'b00000000000000000000000010111011;
					w[216]  = 32'b00000000000000000000000010111000;
					w[217]  = 32'b00000000000000000000000010110101;
					w[218]  = 32'b00000000000000000000000010110010;
					w[219]  = 32'b00000000000000000000000010101111;
					w[220]  = 32'b00000000000000000000000010101100;
					w[221]  = 32'b00000000000000000000000010101000;
					w[222]  = 32'b00000000000000000000000010100101;
					w[223]  = 32'b00000000000000000000000010100010;
					w[224]  = 32'b00000000000000000000000010011111;
					w[225]  = 32'b00000000000000000000000010011100;
					w[226]  = 32'b00000000000000000000000010011001;
					w[227]  = 32'b00000000000000000000000010010101;
					w[228]  = 32'b00000000000000000000000010010010;
					w[229]  = 32'b00000000000000000000000010001111;
					w[230]  = 32'b00000000000000000000000010001100;
					w[231]  = 32'b00000000000000000000000010001001;
					w[232]  = 32'b00000000000000000000000010000101;
					w[233]  = 32'b00000000000000000000000010000010;
					w[234]  = 32'b00000000000000000000000001111111;
					w[235]  = 32'b00000000000000000000000001111100;
					w[236]  = 32'b00000000000000000000000001111001;
					w[237]  = 32'b00000000000000000000000001110101;
					w[238]  = 32'b00000000000000000000000001110010;
					w[239]  = 32'b00000000000000000000000001101111;
					w[240]  = 32'b00000000000000000000000001101100;
					w[241]  = 32'b00000000000000000000000001101001;
					w[242]  = 32'b00000000000000000000000001100110;
					w[243]  = 32'b00000000000000000000000001100011;
					w[244]  = 32'b00000000000000000000000001100000;
					w[245]  = 32'b00000000000000000000000001011101;
					w[246]  = 32'b00000000000000000000000001011010;
					w[247]  = 32'b00000000000000000000000001010111;
					w[248]  = 32'b00000000000000000000000001010100;
					w[249]  = 32'b00000000000000000000000001010001;
					w[250]  = 32'b00000000000000000000000001001110;
					w[251]  = 32'b00000000000000000000000001001011;
					w[252]  = 32'b00000000000000000000000001001000;
					w[253]  = 32'b00000000000000000000000001000101;
					w[254]  = 32'b00000000000000000000000001000011;
					w[255]  = 32'b00000000000000000000000001000000;
					w[256]  = 32'b00000000000000000000000000111101;
					w[257]  = 32'b00000000000000000000000000111011;
					w[258]  = 32'b00000000000000000000000000111000;
					w[259]  = 32'b00000000000000000000000000110110;
					w[260]  = 32'b00000000000000000000000000110011;
					w[261]  = 32'b00000000000000000000000000110001;
					w[262]  = 32'b00000000000000000000000000101110;
					w[263]  = 32'b00000000000000000000000000101100;
					w[264]  = 32'b00000000000000000000000000101010;
					w[265]  = 32'b00000000000000000000000000100111;
					w[266]  = 32'b00000000000000000000000000100101;
					w[267]  = 32'b00000000000000000000000000100011;
					w[268]  = 32'b00000000000000000000000000100001;
					w[269]  = 32'b00000000000000000000000000011111;
					w[270]  = 32'b00000000000000000000000000011101;
					w[271]  = 32'b00000000000000000000000000011011;
					w[272]  = 32'b00000000000000000000000000011001;
					w[273]  = 32'b00000000000000000000000000010111;
					w[274]  = 32'b00000000000000000000000000010110;
					w[275]  = 32'b00000000000000000000000000010100;
					w[276]  = 32'b00000000000000000000000000010010;
					w[277]  = 32'b00000000000000000000000000010001;
					w[278]  = 32'b00000000000000000000000000001111;
					w[279]  = 32'b00000000000000000000000000001110;
					w[280]  = 32'b00000000000000000000000000001100;
					w[281]  = 32'b00000000000000000000000000001011;
					w[282]  = 32'b00000000000000000000000000001010;
					w[283]  = 32'b00000000000000000000000000001001;
					w[284]  = 32'b00000000000000000000000000001000;
					w[285]  = 32'b00000000000000000000000000000111;
					w[286]  = 32'b00000000000000000000000000000110;
					w[287]  = 32'b00000000000000000000000000000101;
					w[288]  = 32'b00000000000000000000000000000100;
					w[289]  = 32'b00000000000000000000000000000011;
					w[290]  = 32'b00000000000000000000000000000010;
					w[291]  = 32'b00000000000000000000000000000010;
					w[292]  = 32'b00000000000000000000000000000001;
					w[293]  = 32'b00000000000000000000000000000001;
					w[294]  = 32'b00000000000000000000000000000000;
					w[295]  = 32'b00000000000000000000000000000000;
					w[296]  = 32'b00000000000000000000000000000000;
					w[297]  = 32'b00000000000000000000000000000000;
					w[298]  = 32'b00000000000000000000000000000000;
					w[299]  = 32'b00000000000000000000000000000000;
					w[300]  = 32'b00000000000000000000000000000000;
					w[301]  = 32'b00000000000000000000000000000000;
					w[302]  = 32'b00000000000000000000000000000000;
					w[303]  = 32'b00000000000000000000000000000000;
					w[304]  = 32'b00000000000000000000000000000000;
					w[305]  = 32'b00000000000000000000000000000000;
					w[306]  = 32'b00000000000000000000000000000000;
					w[307]  = 32'b00000000000000000000000000000000;
					w[308]  = 32'b00000000000000000000000000000000;
					w[309]  = 32'b00000000000000000000000000000000;
					w[310]  = 32'b00000000000000000000000000000000;
					w[311]  = 32'b00000000000000000000000000000000;
					w[312]  = 32'b00000000000000000000000000000000;
					w[313]  = 32'b00000000000000000000000000000000;
					w[314]  = 32'b00000000000000000000000000000000;
					w[315]  = 32'b00000000000000000000000000000000;
					w[316]  = 32'b00000000000000000000000000000000;
					w[317]  = 32'b00000000000000000000000000000000;
					w[318]  = 32'b00000000000000000000000000000000;
					w[319]  = 32'b00000000000000000000000000000000;
	
	
	
		dataout = w[addr];
	end
endmodule
