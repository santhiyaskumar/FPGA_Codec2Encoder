/*
* Module         - ROM_cb3
* Top module     - cbselect
* Project        - CODEC2_ENCODE_2400
* Developer      - Santhiya S
* Date           - Mon Feb 04 15:19:31 2019
*
* Description    -
* Inputs         -
*static const float codes3[] = {
  700,
  800,
  900,
  1000,
  1100,
  1200,
  1300,
  1400,
  1500,
  1600,
  1700,
  1800,
  1900,
  2000,
  2100,
  2200
*};
*32 bits fixed point representation
   S - E  - M
   1 - 15 - 16
*/
module ROM_cb3(addr,dataout);

	parameter N = 32;
	input [3:0] addr;
	output reg [N-1:0] dataout;

	reg [N-1:0] cb3[15:0];
	
	always@(*)
	begin
			cb3[0] = 32'b00000010101111000000000000000000;
			cb3[1] = 32'b00000011001000000000000000000000;
			cb3[2] = 32'b00000011100001000000000000000000;
			cb3[3] = 32'b00000011111010000000000000000000;
			cb3[4] = 32'b00000100010011000000000000000000;
			cb3[5] = 32'b00000100101100000000000000000000;
			cb3[6] = 32'b00000101000101000000000000000000;
			cb3[7] = 32'b00000101011110000000000000000000;
			cb3[8] = 32'b00000101110111000000000000000000;
			cb3[9] = 32'b00000110010000000000000000000000;
			cb3[10] = 32'b00000110101001000000000000000000;
			cb3[11] = 32'b00000111000010000000000000000000;
			cb3[12] = 32'b00000111011011000000000000000000;
			cb3[13] = 32'b00000111110100000000000000000000;
			cb3[14] = 32'b00001000001101000000000000000000;
			cb3[15] = 32'b00001000100110000000000000000000;

		dataout = cb3[addr];
	end
endmodule
